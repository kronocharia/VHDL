
PACKAGE ex4_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
        swapxy,negx,negy: INTEGER; -- swap inputs for octant
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 8000, 8000, 0, 0, 1, 1),
		(start, 8000, 8000, 0, 0, 0, 0, 1, 1),
		(drawing, 8000, 8000, 0, 0, 0, 0, 1, 1),
		(drawing, 7999, 7999, 0, 0, 0, 0, 1, 1),
		(drawing, 7998, 7998, 0, 0, 0, 0, 1, 1),
		(drawing, 7997, 7997, 0, 0, 0, 0, 1, 1),
		(drawing, 7996, 7996, 0, 0, 0, 0, 1, 1),
		(drawing, 7995, 7995, 0, 0, 0, 0, 1, 1),
		(drawing, 7994, 7994, 0, 0, 0, 0, 1, 1),
		(drawing, 7993, 7993, 0, 0, 0, 0, 1, 1),
		(drawing, 7992, 7992, 0, 0, 0, 0, 1, 1),
		(drawing, 7991, 7991, 0, 0, 0, 0, 1, 1),
		(drawing, 7990, 7990, 0, 0, 0, 0, 1, 1),
		(drawing, 7989, 7989, 0, 0, 0, 0, 1, 1),
		(drawing, 7988, 7988, 0, 0, 0, 0, 1, 1),
		(drawing, 7987, 7987, 0, 0, 0, 0, 1, 1),
		(drawing, 7986, 7986, 0, 0, 0, 0, 1, 1),
		(drawing, 7985, 7985, 0, 0, 0, 0, 1, 1),
		(drawing, 7984, 7984, 0, 0, 0, 0, 1, 1),
		(drawing, 7983, 7983, 0, 0, 0, 0, 1, 1),
		(drawing, 7982, 7982, 0, 0, 0, 0, 1, 1),
		(drawing, 7981, 7981, 0, 0, 0, 0, 1, 1),
		(drawing, 7980, 7980, 0, 0, 0, 0, 1, 1),
		(drawing, 7979, 7979, 0, 0, 0, 0, 1, 1),
		(drawing, 7978, 7978, 0, 0, 0, 0, 1, 1),
		(drawing, 7977, 7977, 0, 0, 0, 0, 1, 1),
		(drawing, 7976, 7976, 0, 0, 0, 0, 1, 1),
		(drawing, 7975, 7975, 0, 0, 0, 0, 1, 1),
		(drawing, 7974, 7974, 0, 0, 0, 0, 1, 1),
		(drawing, 7973, 7973, 0, 0, 0, 0, 1, 1),
		(drawing, 7972, 7972, 0, 0, 0, 0, 1, 1),
		(drawing, 7971, 7971, 0, 0, 0, 0, 1, 1),
		(drawing, 7970, 7970, 0, 0, 0, 0, 1, 1),
		(drawing, 7969, 7969, 0, 0, 0, 0, 1, 1),
		(drawing, 7968, 7968, 0, 0, 0, 0, 1, 1),
		(drawing, 7967, 7967, 0, 0, 0, 0, 1, 1),
		(drawing, 7966, 7966, 0, 0, 0, 0, 1, 1),
		(drawing, 7965, 7965, 0, 0, 0, 0, 1, 1),
		(drawing, 7964, 7964, 0, 0, 0, 0, 1, 1),
		(drawing, 7963, 7963, 0, 0, 0, 0, 1, 1),
		(drawing, 7962, 7962, 0, 0, 0, 0, 1, 1),
		(drawing, 7961, 7961, 0, 0, 0, 0, 1, 1),
		(drawing, 7960, 7960, 0, 0, 0, 0, 1, 1),
		(drawing, 7959, 7959, 0, 0, 0, 0, 1, 1),
		(drawing, 7958, 7958, 0, 0, 0, 0, 1, 1),
		(drawing, 7957, 7957, 0, 0, 0, 0, 1, 1),
		(drawing, 7956, 7956, 0, 0, 0, 0, 1, 1),
		(drawing, 7955, 7955, 0, 0, 0, 0, 1, 1),
		(drawing, 7954, 7954, 0, 0, 0, 0, 1, 1),
		(drawing, 7953, 7953, 0, 0, 0, 0, 1, 1),
		(drawing, 7952, 7952, 0, 0, 0, 0, 1, 1),
		(drawing, 7951, 7951, 0, 0, 0, 0, 1, 1),
		(drawing, 7950, 7950, 0, 0, 0, 0, 1, 1),
		(drawing, 7949, 7949, 0, 0, 0, 0, 1, 1),
		(drawing, 7948, 7948, 0, 0, 0, 0, 1, 1),
		(drawing, 7947, 7947, 0, 0, 0, 0, 1, 1),
		(drawing, 7946, 7946, 0, 0, 0, 0, 1, 1),
		(drawing, 7945, 7945, 0, 0, 0, 0, 1, 1),
		(drawing, 7944, 7944, 0, 0, 0, 0, 1, 1),
		(drawing, 7943, 7943, 0, 0, 0, 0, 1, 1),
		(drawing, 7942, 7942, 0, 0, 0, 0, 1, 1),
		(drawing, 7941, 7941, 0, 0, 0, 0, 1, 1),
		(drawing, 7940, 7940, 0, 0, 0, 0, 1, 1),
		(drawing, 7939, 7939, 0, 0, 0, 0, 1, 1),
		(drawing, 7938, 7938, 0, 0, 0, 0, 1, 1),
		(drawing, 7937, 7937, 0, 0, 0, 0, 1, 1),
		(drawing, 7936, 7936, 0, 0, 0, 0, 1, 1),
		(drawing, 7935, 7935, 0, 0, 0, 0, 1, 1),
		(drawing, 7934, 7934, 0, 0, 0, 0, 1, 1),
		(drawing, 7933, 7933, 0, 0, 0, 0, 1, 1),
		(drawing, 7932, 7932, 0, 0, 0, 0, 1, 1),
		(drawing, 7931, 7931, 0, 0, 0, 0, 1, 1),
		(drawing, 7930, 7930, 0, 0, 0, 0, 1, 1),
		(drawing, 7929, 7929, 0, 0, 0, 0, 1, 1),
		(drawing, 7928, 7928, 0, 0, 0, 0, 1, 1),
		(drawing, 7927, 7927, 0, 0, 0, 0, 1, 1),
		(drawing, 7926, 7926, 0, 0, 0, 0, 1, 1),
		(drawing, 7925, 7925, 0, 0, 0, 0, 1, 1),
		(drawing, 7924, 7924, 0, 0, 0, 0, 1, 1),
		(drawing, 7923, 7923, 0, 0, 0, 0, 1, 1),
		(drawing, 7922, 7922, 0, 0, 0, 0, 1, 1),
		(drawing, 7921, 7921, 0, 0, 0, 0, 1, 1),
		(drawing, 7920, 7920, 0, 0, 0, 0, 1, 1),
		(drawing, 7919, 7919, 0, 0, 0, 0, 1, 1),
		(drawing, 7918, 7918, 0, 0, 0, 0, 1, 1),
		(drawing, 7917, 7917, 0, 0, 0, 0, 1, 1),
		(drawing, 7916, 7916, 0, 0, 0, 0, 1, 1),
		(drawing, 7915, 7915, 0, 0, 0, 0, 1, 1),
		(drawing, 7914, 7914, 0, 0, 0, 0, 1, 1),
		(drawing, 7913, 7913, 0, 0, 0, 0, 1, 1),
		(drawing, 7912, 7912, 0, 0, 0, 0, 1, 1),
		(drawing, 7911, 7911, 0, 0, 0, 0, 1, 1),
		(drawing, 7910, 7910, 0, 0, 0, 0, 1, 1),
		(drawing, 7909, 7909, 0, 0, 0, 0, 1, 1),
		(drawing, 7908, 7908, 0, 0, 0, 0, 1, 1),
		(drawing, 7907, 7907, 0, 0, 0, 0, 1, 1),
		(drawing, 7906, 7906, 0, 0, 0, 0, 1, 1),
		(drawing, 7905, 7905, 0, 0, 0, 0, 1, 1),
		(drawing, 7904, 7904, 0, 0, 0, 0, 1, 1),
		(drawing, 7903, 7903, 0, 0, 0, 0, 1, 1),
		(drawing, 7902, 7902, 0, 0, 0, 0, 1, 1),
		(drawing, 7901, 7901, 0, 0, 0, 0, 1, 1),
		(drawing, 7900, 7900, 0, 0, 0, 0, 1, 1),
		(drawing, 7899, 7899, 0, 0, 0, 0, 1, 1),
		(drawing, 7898, 7898, 0, 0, 0, 0, 1, 1),
		(drawing, 7897, 7897, 0, 0, 0, 0, 1, 1),
		(drawing, 7896, 7896, 0, 0, 0, 0, 1, 1),
		(drawing, 7895, 7895, 0, 0, 0, 0, 1, 1),
		(drawing, 7894, 7894, 0, 0, 0, 0, 1, 1),
		(drawing, 7893, 7893, 0, 0, 0, 0, 1, 1),
		(drawing, 7892, 7892, 0, 0, 0, 0, 1, 1),
		(drawing, 7891, 7891, 0, 0, 0, 0, 1, 1),
		(drawing, 7890, 7890, 0, 0, 0, 0, 1, 1),
		(drawing, 7889, 7889, 0, 0, 0, 0, 1, 1),
		(drawing, 7888, 7888, 0, 0, 0, 0, 1, 1),
		(drawing, 7887, 7887, 0, 0, 0, 0, 1, 1),
		(drawing, 7886, 7886, 0, 0, 0, 0, 1, 1),
		(drawing, 7885, 7885, 0, 0, 0, 0, 1, 1),
		(drawing, 7884, 7884, 0, 0, 0, 0, 1, 1),
		(drawing, 7883, 7883, 0, 0, 0, 0, 1, 1),
		(drawing, 7882, 7882, 0, 0, 0, 0, 1, 1),
		(drawing, 7881, 7881, 0, 0, 0, 0, 1, 1),
		(drawing, 7880, 7880, 0, 0, 0, 0, 1, 1),
		(drawing, 7879, 7879, 0, 0, 0, 0, 1, 1),
		(drawing, 7878, 7878, 0, 0, 0, 0, 1, 1),
		(drawing, 7877, 7877, 0, 0, 0, 0, 1, 1),
		(drawing, 7876, 7876, 0, 0, 0, 0, 1, 1),
		(drawing, 7875, 7875, 0, 0, 0, 0, 1, 1),
		(drawing, 7874, 7874, 0, 0, 0, 0, 1, 1),
		(drawing, 7873, 7873, 0, 0, 0, 0, 1, 1),
		(drawing, 7872, 7872, 0, 0, 0, 0, 1, 1),
		(drawing, 7871, 7871, 0, 0, 0, 0, 1, 1),
		(drawing, 7870, 7870, 0, 0, 0, 0, 1, 1),
		(drawing, 7869, 7869, 0, 0, 0, 0, 1, 1),
		(drawing, 7868, 7868, 0, 0, 0, 0, 1, 1),
		(drawing, 7867, 7867, 0, 0, 0, 0, 1, 1),
		(drawing, 7866, 7866, 0, 0, 0, 0, 1, 1),
		(drawing, 7865, 7865, 0, 0, 0, 0, 1, 1),
		(drawing, 7864, 7864, 0, 0, 0, 0, 1, 1),
		(drawing, 7863, 7863, 0, 0, 0, 0, 1, 1),
		(drawing, 7862, 7862, 0, 0, 0, 0, 1, 1),
		(drawing, 7861, 7861, 0, 0, 0, 0, 1, 1),
		(drawing, 7860, 7860, 0, 0, 0, 0, 1, 1),
		(drawing, 7859, 7859, 0, 0, 0, 0, 1, 1),
		(drawing, 7858, 7858, 0, 0, 0, 0, 1, 1),
		(drawing, 7857, 7857, 0, 0, 0, 0, 1, 1),
		(drawing, 7856, 7856, 0, 0, 0, 0, 1, 1),
		(drawing, 7855, 7855, 0, 0, 0, 0, 1, 1),
		(drawing, 7854, 7854, 0, 0, 0, 0, 1, 1),
		(drawing, 7853, 7853, 0, 0, 0, 0, 1, 1),
		(drawing, 7852, 7852, 0, 0, 0, 0, 1, 1),
		(drawing, 7851, 7851, 0, 0, 0, 0, 1, 1),
		(drawing, 7850, 7850, 0, 0, 0, 0, 1, 1),
		(drawing, 7849, 7849, 0, 0, 0, 0, 1, 1),
		(drawing, 7848, 7848, 0, 0, 0, 0, 1, 1),
		(drawing, 7847, 7847, 0, 0, 0, 0, 1, 1),
		(drawing, 7846, 7846, 0, 0, 0, 0, 1, 1),
		(drawing, 7845, 7845, 0, 0, 0, 0, 1, 1),
		(drawing, 7844, 7844, 0, 0, 0, 0, 1, 1),
		(drawing, 7843, 7843, 0, 0, 0, 0, 1, 1),
		(drawing, 7842, 7842, 0, 0, 0, 0, 1, 1),
		(drawing, 7841, 7841, 0, 0, 0, 0, 1, 1),
		(drawing, 7840, 7840, 0, 0, 0, 0, 1, 1),
		(drawing, 7839, 7839, 0, 0, 0, 0, 1, 1),
		(drawing, 7838, 7838, 0, 0, 0, 0, 1, 1),
		(drawing, 7837, 7837, 0, 0, 0, 0, 1, 1),
		(drawing, 7836, 7836, 0, 0, 0, 0, 1, 1),
		(drawing, 7835, 7835, 0, 0, 0, 0, 1, 1),
		(drawing, 7834, 7834, 0, 0, 0, 0, 1, 1),
		(drawing, 7833, 7833, 0, 0, 0, 0, 1, 1),
		(drawing, 7832, 7832, 0, 0, 0, 0, 1, 1),
		(drawing, 7831, 7831, 0, 0, 0, 0, 1, 1),
		(drawing, 7830, 7830, 0, 0, 0, 0, 1, 1),
		(drawing, 7829, 7829, 0, 0, 0, 0, 1, 1),
		(drawing, 7828, 7828, 0, 0, 0, 0, 1, 1),
		(drawing, 7827, 7827, 0, 0, 0, 0, 1, 1),
		(drawing, 7826, 7826, 0, 0, 0, 0, 1, 1),
		(drawing, 7825, 7825, 0, 0, 0, 0, 1, 1),
		(drawing, 7824, 7824, 0, 0, 0, 0, 1, 1),
		(drawing, 7823, 7823, 0, 0, 0, 0, 1, 1),
		(drawing, 7822, 7822, 0, 0, 0, 0, 1, 1),
		(drawing, 7821, 7821, 0, 0, 0, 0, 1, 1),
		(drawing, 7820, 7820, 0, 0, 0, 0, 1, 1),
		(drawing, 7819, 7819, 0, 0, 0, 0, 1, 1),
		(drawing, 7818, 7818, 0, 0, 0, 0, 1, 1),
		(drawing, 7817, 7817, 0, 0, 0, 0, 1, 1),
		(drawing, 7816, 7816, 0, 0, 0, 0, 1, 1),
		(drawing, 7815, 7815, 0, 0, 0, 0, 1, 1),
		(drawing, 7814, 7814, 0, 0, 0, 0, 1, 1),
		(drawing, 7813, 7813, 0, 0, 0, 0, 1, 1),
		(drawing, 7812, 7812, 0, 0, 0, 0, 1, 1),
		(drawing, 7811, 7811, 0, 0, 0, 0, 1, 1),
		(drawing, 7810, 7810, 0, 0, 0, 0, 1, 1),
		(drawing, 7809, 7809, 0, 0, 0, 0, 1, 1),
		(drawing, 7808, 7808, 0, 0, 0, 0, 1, 1),
		(drawing, 7807, 7807, 0, 0, 0, 0, 1, 1),
		(drawing, 7806, 7806, 0, 0, 0, 0, 1, 1),
		(drawing, 7805, 7805, 0, 0, 0, 0, 1, 1),
		(drawing, 7804, 7804, 0, 0, 0, 0, 1, 1),
		(drawing, 7803, 7803, 0, 0, 0, 0, 1, 1),
		(drawing, 7802, 7802, 0, 0, 0, 0, 1, 1),
		(drawing, 7801, 7801, 0, 0, 0, 0, 1, 1),
		(drawing, 7800, 7800, 0, 0, 0, 0, 1, 1),
		(drawing, 7799, 7799, 0, 0, 0, 0, 1, 1),
		(drawing, 7798, 7798, 0, 0, 0, 0, 1, 1),
		(drawing, 7797, 7797, 0, 0, 0, 0, 1, 1),
		(drawing, 7796, 7796, 0, 0, 0, 0, 1, 1),
		(drawing, 7795, 7795, 0, 0, 0, 0, 1, 1),
		(drawing, 7794, 7794, 0, 0, 0, 0, 1, 1),
		(drawing, 7793, 7793, 0, 0, 0, 0, 1, 1),
		(drawing, 7792, 7792, 0, 0, 0, 0, 1, 1),
		(drawing, 7791, 7791, 0, 0, 0, 0, 1, 1),
		(drawing, 7790, 7790, 0, 0, 0, 0, 1, 1),
		(drawing, 7789, 7789, 0, 0, 0, 0, 1, 1),
		(drawing, 7788, 7788, 0, 0, 0, 0, 1, 1),
		(drawing, 7787, 7787, 0, 0, 0, 0, 1, 1),
		(drawing, 7786, 7786, 0, 0, 0, 0, 1, 1),
		(drawing, 7785, 7785, 0, 0, 0, 0, 1, 1),
		(drawing, 7784, 7784, 0, 0, 0, 0, 1, 1),
		(drawing, 7783, 7783, 0, 0, 0, 0, 1, 1),
		(drawing, 7782, 7782, 0, 0, 0, 0, 1, 1),
		(drawing, 7781, 7781, 0, 0, 0, 0, 1, 1),
		(drawing, 7780, 7780, 0, 0, 0, 0, 1, 1),
		(drawing, 7779, 7779, 0, 0, 0, 0, 1, 1),
		(drawing, 7778, 7778, 0, 0, 0, 0, 1, 1),
		(drawing, 7777, 7777, 0, 0, 0, 0, 1, 1),
		(drawing, 7776, 7776, 0, 0, 0, 0, 1, 1),
		(drawing, 7775, 7775, 0, 0, 0, 0, 1, 1),
		(drawing, 7774, 7774, 0, 0, 0, 0, 1, 1),
		(drawing, 7773, 7773, 0, 0, 0, 0, 1, 1),
		(drawing, 7772, 7772, 0, 0, 0, 0, 1, 1),
		(drawing, 7771, 7771, 0, 0, 0, 0, 1, 1),
		(drawing, 7770, 7770, 0, 0, 0, 0, 1, 1),
		(drawing, 7769, 7769, 0, 0, 0, 0, 1, 1),
		(drawing, 7768, 7768, 0, 0, 0, 0, 1, 1),
		(drawing, 7767, 7767, 0, 0, 0, 0, 1, 1),
		(drawing, 7766, 7766, 0, 0, 0, 0, 1, 1),
		(drawing, 7765, 7765, 0, 0, 0, 0, 1, 1),
		(drawing, 7764, 7764, 0, 0, 0, 0, 1, 1),
		(drawing, 7763, 7763, 0, 0, 0, 0, 1, 1),
		(drawing, 7762, 7762, 0, 0, 0, 0, 1, 1),
		(drawing, 7761, 7761, 0, 0, 0, 0, 1, 1),
		(drawing, 7760, 7760, 0, 0, 0, 0, 1, 1),
		(drawing, 7759, 7759, 0, 0, 0, 0, 1, 1),
		(drawing, 7758, 7758, 0, 0, 0, 0, 1, 1),
		(drawing, 7757, 7757, 0, 0, 0, 0, 1, 1),
		(drawing, 7756, 7756, 0, 0, 0, 0, 1, 1),
		(drawing, 7755, 7755, 0, 0, 0, 0, 1, 1),
		(drawing, 7754, 7754, 0, 0, 0, 0, 1, 1),
		(drawing, 7753, 7753, 0, 0, 0, 0, 1, 1),
		(drawing, 7752, 7752, 0, 0, 0, 0, 1, 1),
		(drawing, 7751, 7751, 0, 0, 0, 0, 1, 1),
		(drawing, 7750, 7750, 0, 0, 0, 0, 1, 1),
		(drawing, 7749, 7749, 0, 0, 0, 0, 1, 1),
		(drawing, 7748, 7748, 0, 0, 0, 0, 1, 1),
		(drawing, 7747, 7747, 0, 0, 0, 0, 1, 1),
		(drawing, 7746, 7746, 0, 0, 0, 0, 1, 1),
		(drawing, 7745, 7745, 0, 0, 0, 0, 1, 1),
		(drawing, 7744, 7744, 0, 0, 0, 0, 1, 1),
		(drawing, 7743, 7743, 0, 0, 0, 0, 1, 1),
		(drawing, 7742, 7742, 0, 0, 0, 0, 1, 1),
		(drawing, 7741, 7741, 0, 0, 0, 0, 1, 1),
		(drawing, 7740, 7740, 0, 0, 0, 0, 1, 1),
		(drawing, 7739, 7739, 0, 0, 0, 0, 1, 1),
		(drawing, 7738, 7738, 0, 0, 0, 0, 1, 1),
		(drawing, 7737, 7737, 0, 0, 0, 0, 1, 1),
		(drawing, 7736, 7736, 0, 0, 0, 0, 1, 1),
		(drawing, 7735, 7735, 0, 0, 0, 0, 1, 1),
		(drawing, 7734, 7734, 0, 0, 0, 0, 1, 1),
		(drawing, 7733, 7733, 0, 0, 0, 0, 1, 1),
		(drawing, 7732, 7732, 0, 0, 0, 0, 1, 1),
		(drawing, 7731, 7731, 0, 0, 0, 0, 1, 1),
		(drawing, 7730, 7730, 0, 0, 0, 0, 1, 1),
		(drawing, 7729, 7729, 0, 0, 0, 0, 1, 1),
		(drawing, 7728, 7728, 0, 0, 0, 0, 1, 1),
		(drawing, 7727, 7727, 0, 0, 0, 0, 1, 1),
		(drawing, 7726, 7726, 0, 0, 0, 0, 1, 1),
		(drawing, 7725, 7725, 0, 0, 0, 0, 1, 1),
		(drawing, 7724, 7724, 0, 0, 0, 0, 1, 1),
		(drawing, 7723, 7723, 0, 0, 0, 0, 1, 1),
		(drawing, 7722, 7722, 0, 0, 0, 0, 1, 1),
		(drawing, 7721, 7721, 0, 0, 0, 0, 1, 1),
		(drawing, 7720, 7720, 0, 0, 0, 0, 1, 1),
		(drawing, 7719, 7719, 0, 0, 0, 0, 1, 1),
		(drawing, 7718, 7718, 0, 0, 0, 0, 1, 1),
		(drawing, 7717, 7717, 0, 0, 0, 0, 1, 1),
		(drawing, 7716, 7716, 0, 0, 0, 0, 1, 1),
		(drawing, 7715, 7715, 0, 0, 0, 0, 1, 1),
		(drawing, 7714, 7714, 0, 0, 0, 0, 1, 1),
		(drawing, 7713, 7713, 0, 0, 0, 0, 1, 1),
		(drawing, 7712, 7712, 0, 0, 0, 0, 1, 1),
		(drawing, 7711, 7711, 0, 0, 0, 0, 1, 1),
		(drawing, 7710, 7710, 0, 0, 0, 0, 1, 1),
		(drawing, 7709, 7709, 0, 0, 0, 0, 1, 1),
		(drawing, 7708, 7708, 0, 0, 0, 0, 1, 1),
		(drawing, 7707, 7707, 0, 0, 0, 0, 1, 1),
		(drawing, 7706, 7706, 0, 0, 0, 0, 1, 1),
		(drawing, 7705, 7705, 0, 0, 0, 0, 1, 1),
		(drawing, 7704, 7704, 0, 0, 0, 0, 1, 1),
		(drawing, 7703, 7703, 0, 0, 0, 0, 1, 1),
		(drawing, 7702, 7702, 0, 0, 0, 0, 1, 1),
		(drawing, 7701, 7701, 0, 0, 0, 0, 1, 1),
		(drawing, 7700, 7700, 0, 0, 0, 0, 1, 1),
		(drawing, 7699, 7699, 0, 0, 0, 0, 1, 1),
		(drawing, 7698, 7698, 0, 0, 0, 0, 1, 1),
		(drawing, 7697, 7697, 0, 0, 0, 0, 1, 1),
		(drawing, 7696, 7696, 0, 0, 0, 0, 1, 1),
		(drawing, 7695, 7695, 0, 0, 0, 0, 1, 1),
		(drawing, 7694, 7694, 0, 0, 0, 0, 1, 1),
		(drawing, 7693, 7693, 0, 0, 0, 0, 1, 1),
		(drawing, 7692, 7692, 0, 0, 0, 0, 1, 1),
		(drawing, 7691, 7691, 0, 0, 0, 0, 1, 1),
		(drawing, 7690, 7690, 0, 0, 0, 0, 1, 1),
		(drawing, 7689, 7689, 0, 0, 0, 0, 1, 1),
		(drawing, 7688, 7688, 0, 0, 0, 0, 1, 1),
		(drawing, 7687, 7687, 0, 0, 0, 0, 1, 1),
		(drawing, 7686, 7686, 0, 0, 0, 0, 1, 1),
		(drawing, 7685, 7685, 0, 0, 0, 0, 1, 1),
		(drawing, 7684, 7684, 0, 0, 0, 0, 1, 1),
		(drawing, 7683, 7683, 0, 0, 0, 0, 1, 1),
		(drawing, 7682, 7682, 0, 0, 0, 0, 1, 1),
		(drawing, 7681, 7681, 0, 0, 0, 0, 1, 1),
		(drawing, 7680, 7680, 0, 0, 0, 0, 1, 1),
		(drawing, 7679, 7679, 0, 0, 0, 0, 1, 1),
		(drawing, 7678, 7678, 0, 0, 0, 0, 1, 1),
		(drawing, 7677, 7677, 0, 0, 0, 0, 1, 1),
		(drawing, 7676, 7676, 0, 0, 0, 0, 1, 1),
		(drawing, 7675, 7675, 0, 0, 0, 0, 1, 1),
		(drawing, 7674, 7674, 0, 0, 0, 0, 1, 1),
		(drawing, 7673, 7673, 0, 0, 0, 0, 1, 1),
		(drawing, 7672, 7672, 0, 0, 0, 0, 1, 1),
		(drawing, 7671, 7671, 0, 0, 0, 0, 1, 1),
		(drawing, 7670, 7670, 0, 0, 0, 0, 1, 1),
		(drawing, 7669, 7669, 0, 0, 0, 0, 1, 1),
		(drawing, 7668, 7668, 0, 0, 0, 0, 1, 1),
		(drawing, 7667, 7667, 0, 0, 0, 0, 1, 1),
		(drawing, 7666, 7666, 0, 0, 0, 0, 1, 1),
		(drawing, 7665, 7665, 0, 0, 0, 0, 1, 1),
		(drawing, 7664, 7664, 0, 0, 0, 0, 1, 1),
		(drawing, 7663, 7663, 0, 0, 0, 0, 1, 1),
		(drawing, 7662, 7662, 0, 0, 0, 0, 1, 1),
		(drawing, 7661, 7661, 0, 0, 0, 0, 1, 1),
		(drawing, 7660, 7660, 0, 0, 0, 0, 1, 1),
		(drawing, 7659, 7659, 0, 0, 0, 0, 1, 1),
		(drawing, 7658, 7658, 0, 0, 0, 0, 1, 1),
		(drawing, 7657, 7657, 0, 0, 0, 0, 1, 1),
		(drawing, 7656, 7656, 0, 0, 0, 0, 1, 1),
		(drawing, 7655, 7655, 0, 0, 0, 0, 1, 1),
		(drawing, 7654, 7654, 0, 0, 0, 0, 1, 1),
		(drawing, 7653, 7653, 0, 0, 0, 0, 1, 1),
		(drawing, 7652, 7652, 0, 0, 0, 0, 1, 1),
		(drawing, 7651, 7651, 0, 0, 0, 0, 1, 1),
		(drawing, 7650, 7650, 0, 0, 0, 0, 1, 1),
		(drawing, 7649, 7649, 0, 0, 0, 0, 1, 1),
		(drawing, 7648, 7648, 0, 0, 0, 0, 1, 1),
		(drawing, 7647, 7647, 0, 0, 0, 0, 1, 1),
		(drawing, 7646, 7646, 0, 0, 0, 0, 1, 1),
		(drawing, 7645, 7645, 0, 0, 0, 0, 1, 1),
		(drawing, 7644, 7644, 0, 0, 0, 0, 1, 1),
		(drawing, 7643, 7643, 0, 0, 0, 0, 1, 1),
		(drawing, 7642, 7642, 0, 0, 0, 0, 1, 1),
		(drawing, 7641, 7641, 0, 0, 0, 0, 1, 1),
		(drawing, 7640, 7640, 0, 0, 0, 0, 1, 1),
		(drawing, 7639, 7639, 0, 0, 0, 0, 1, 1),
		(drawing, 7638, 7638, 0, 0, 0, 0, 1, 1),
		(drawing, 7637, 7637, 0, 0, 0, 0, 1, 1),
		(drawing, 7636, 7636, 0, 0, 0, 0, 1, 1),
		(drawing, 7635, 7635, 0, 0, 0, 0, 1, 1),
		(drawing, 7634, 7634, 0, 0, 0, 0, 1, 1),
		(drawing, 7633, 7633, 0, 0, 0, 0, 1, 1),
		(drawing, 7632, 7632, 0, 0, 0, 0, 1, 1),
		(drawing, 7631, 7631, 0, 0, 0, 0, 1, 1),
		(drawing, 7630, 7630, 0, 0, 0, 0, 1, 1),
		(drawing, 7629, 7629, 0, 0, 0, 0, 1, 1),
		(drawing, 7628, 7628, 0, 0, 0, 0, 1, 1),
		(drawing, 7627, 7627, 0, 0, 0, 0, 1, 1),
		(drawing, 7626, 7626, 0, 0, 0, 0, 1, 1),
		(drawing, 7625, 7625, 0, 0, 0, 0, 1, 1),
		(drawing, 7624, 7624, 0, 0, 0, 0, 1, 1),
		(drawing, 7623, 7623, 0, 0, 0, 0, 1, 1),
		(drawing, 7622, 7622, 0, 0, 0, 0, 1, 1),
		(drawing, 7621, 7621, 0, 0, 0, 0, 1, 1),
		(drawing, 7620, 7620, 0, 0, 0, 0, 1, 1),
		(drawing, 7619, 7619, 0, 0, 0, 0, 1, 1),
		(drawing, 7618, 7618, 0, 0, 0, 0, 1, 1),
		(drawing, 7617, 7617, 0, 0, 0, 0, 1, 1),
		(drawing, 7616, 7616, 0, 0, 0, 0, 1, 1),
		(drawing, 7615, 7615, 0, 0, 0, 0, 1, 1),
		(drawing, 7614, 7614, 0, 0, 0, 0, 1, 1),
		(drawing, 7613, 7613, 0, 0, 0, 0, 1, 1),
		(drawing, 7612, 7612, 0, 0, 0, 0, 1, 1),
		(drawing, 7611, 7611, 0, 0, 0, 0, 1, 1),
		(drawing, 7610, 7610, 0, 0, 0, 0, 1, 1),
		(drawing, 7609, 7609, 0, 0, 0, 0, 1, 1),
		(drawing, 7608, 7608, 0, 0, 0, 0, 1, 1),
		(drawing, 7607, 7607, 0, 0, 0, 0, 1, 1),
		(drawing, 7606, 7606, 0, 0, 0, 0, 1, 1),
		(drawing, 7605, 7605, 0, 0, 0, 0, 1, 1),
		(drawing, 7604, 7604, 0, 0, 0, 0, 1, 1),
		(drawing, 7603, 7603, 0, 0, 0, 0, 1, 1),
		(drawing, 7602, 7602, 0, 0, 0, 0, 1, 1),
		(drawing, 7601, 7601, 0, 0, 0, 0, 1, 1),
		(drawing, 7600, 7600, 0, 0, 0, 0, 1, 1),
		(drawing, 7599, 7599, 0, 0, 0, 0, 1, 1),
		(drawing, 7598, 7598, 0, 0, 0, 0, 1, 1),
		(drawing, 7597, 7597, 0, 0, 0, 0, 1, 1),
		(drawing, 7596, 7596, 0, 0, 0, 0, 1, 1),
		(drawing, 7595, 7595, 0, 0, 0, 0, 1, 1),
		(drawing, 7594, 7594, 0, 0, 0, 0, 1, 1),
		(drawing, 7593, 7593, 0, 0, 0, 0, 1, 1),
		(drawing, 7592, 7592, 0, 0, 0, 0, 1, 1),
		(drawing, 7591, 7591, 0, 0, 0, 0, 1, 1),
		(drawing, 7590, 7590, 0, 0, 0, 0, 1, 1),
		(drawing, 7589, 7589, 0, 0, 0, 0, 1, 1),
		(drawing, 7588, 7588, 0, 0, 0, 0, 1, 1),
		(drawing, 7587, 7587, 0, 0, 0, 0, 1, 1),
		(drawing, 7586, 7586, 0, 0, 0, 0, 1, 1),
		(drawing, 7585, 7585, 0, 0, 0, 0, 1, 1),
		(drawing, 7584, 7584, 0, 0, 0, 0, 1, 1),
		(drawing, 7583, 7583, 0, 0, 0, 0, 1, 1),
		(drawing, 7582, 7582, 0, 0, 0, 0, 1, 1),
		(drawing, 7581, 7581, 0, 0, 0, 0, 1, 1),
		(drawing, 7580, 7580, 0, 0, 0, 0, 1, 1),
		(drawing, 7579, 7579, 0, 0, 0, 0, 1, 1),
		(drawing, 7578, 7578, 0, 0, 0, 0, 1, 1),
		(drawing, 7577, 7577, 0, 0, 0, 0, 1, 1),
		(drawing, 7576, 7576, 0, 0, 0, 0, 1, 1),
		(drawing, 7575, 7575, 0, 0, 0, 0, 1, 1),
		(drawing, 7574, 7574, 0, 0, 0, 0, 1, 1),
		(drawing, 7573, 7573, 0, 0, 0, 0, 1, 1),
		(drawing, 7572, 7572, 0, 0, 0, 0, 1, 1),
		(drawing, 7571, 7571, 0, 0, 0, 0, 1, 1),
		(drawing, 7570, 7570, 0, 0, 0, 0, 1, 1),
		(drawing, 7569, 7569, 0, 0, 0, 0, 1, 1),
		(drawing, 7568, 7568, 0, 0, 0, 0, 1, 1),
		(drawing, 7567, 7567, 0, 0, 0, 0, 1, 1),
		(drawing, 7566, 7566, 0, 0, 0, 0, 1, 1),
		(drawing, 7565, 7565, 0, 0, 0, 0, 1, 1),
		(drawing, 7564, 7564, 0, 0, 0, 0, 1, 1),
		(drawing, 7563, 7563, 0, 0, 0, 0, 1, 1),
		(drawing, 7562, 7562, 0, 0, 0, 0, 1, 1),
		(drawing, 7561, 7561, 0, 0, 0, 0, 1, 1),
		(drawing, 7560, 7560, 0, 0, 0, 0, 1, 1),
		(drawing, 7559, 7559, 0, 0, 0, 0, 1, 1),
		(drawing, 7558, 7558, 0, 0, 0, 0, 1, 1),
		(drawing, 7557, 7557, 0, 0, 0, 0, 1, 1),
		(drawing, 7556, 7556, 0, 0, 0, 0, 1, 1),
		(drawing, 7555, 7555, 0, 0, 0, 0, 1, 1),
		(drawing, 7554, 7554, 0, 0, 0, 0, 1, 1),
		(drawing, 7553, 7553, 0, 0, 0, 0, 1, 1),
		(drawing, 7552, 7552, 0, 0, 0, 0, 1, 1),
		(drawing, 7551, 7551, 0, 0, 0, 0, 1, 1),
		(drawing, 7550, 7550, 0, 0, 0, 0, 1, 1),
		(drawing, 7549, 7549, 0, 0, 0, 0, 1, 1),
		(drawing, 7548, 7548, 0, 0, 0, 0, 1, 1),
		(drawing, 7547, 7547, 0, 0, 0, 0, 1, 1),
		(drawing, 7546, 7546, 0, 0, 0, 0, 1, 1),
		(drawing, 7545, 7545, 0, 0, 0, 0, 1, 1),
		(drawing, 7544, 7544, 0, 0, 0, 0, 1, 1),
		(drawing, 7543, 7543, 0, 0, 0, 0, 1, 1),
		(drawing, 7542, 7542, 0, 0, 0, 0, 1, 1),
		(drawing, 7541, 7541, 0, 0, 0, 0, 1, 1),
		(drawing, 7540, 7540, 0, 0, 0, 0, 1, 1),
		(drawing, 7539, 7539, 0, 0, 0, 0, 1, 1),
		(drawing, 7538, 7538, 0, 0, 0, 0, 1, 1),
		(drawing, 7537, 7537, 0, 0, 0, 0, 1, 1),
		(drawing, 7536, 7536, 0, 0, 0, 0, 1, 1),
		(drawing, 7535, 7535, 0, 0, 0, 0, 1, 1),
		(drawing, 7534, 7534, 0, 0, 0, 0, 1, 1),
		(drawing, 7533, 7533, 0, 0, 0, 0, 1, 1),
		(drawing, 7532, 7532, 0, 0, 0, 0, 1, 1),
		(drawing, 7531, 7531, 0, 0, 0, 0, 1, 1),
		(drawing, 7530, 7530, 0, 0, 0, 0, 1, 1),
		(drawing, 7529, 7529, 0, 0, 0, 0, 1, 1),
		(drawing, 7528, 7528, 0, 0, 0, 0, 1, 1),
		(drawing, 7527, 7527, 0, 0, 0, 0, 1, 1),
		(drawing, 7526, 7526, 0, 0, 0, 0, 1, 1),
		(drawing, 7525, 7525, 0, 0, 0, 0, 1, 1),
		(drawing, 7524, 7524, 0, 0, 0, 0, 1, 1),
		(drawing, 7523, 7523, 0, 0, 0, 0, 1, 1),
		(drawing, 7522, 7522, 0, 0, 0, 0, 1, 1),
		(drawing, 7521, 7521, 0, 0, 0, 0, 1, 1),
		(drawing, 7520, 7520, 0, 0, 0, 0, 1, 1),
		(drawing, 7519, 7519, 0, 0, 0, 0, 1, 1),
		(drawing, 7518, 7518, 0, 0, 0, 0, 1, 1),
		(drawing, 7517, 7517, 0, 0, 0, 0, 1, 1),
		(drawing, 7516, 7516, 0, 0, 0, 0, 1, 1),
		(drawing, 7515, 7515, 0, 0, 0, 0, 1, 1),
		(drawing, 7514, 7514, 0, 0, 0, 0, 1, 1),
		(drawing, 7513, 7513, 0, 0, 0, 0, 1, 1),
		(drawing, 7512, 7512, 0, 0, 0, 0, 1, 1),
		(drawing, 7511, 7511, 0, 0, 0, 0, 1, 1),
		(drawing, 7510, 7510, 0, 0, 0, 0, 1, 1),
		(drawing, 7509, 7509, 0, 0, 0, 0, 1, 1),
		(drawing, 7508, 7508, 0, 0, 0, 0, 1, 1),
		(drawing, 7507, 7507, 0, 0, 0, 0, 1, 1),
		(drawing, 7506, 7506, 0, 0, 0, 0, 1, 1),
		(drawing, 7505, 7505, 0, 0, 0, 0, 1, 1),
		(drawing, 7504, 7504, 0, 0, 0, 0, 1, 1),
		(drawing, 7503, 7503, 0, 0, 0, 0, 1, 1),
		(drawing, 7502, 7502, 0, 0, 0, 0, 1, 1),
		(drawing, 7501, 7501, 0, 0, 0, 0, 1, 1),
		(drawing, 7500, 7500, 0, 0, 0, 0, 1, 1),
		(drawing, 7499, 7499, 0, 0, 0, 0, 1, 1),
		(drawing, 7498, 7498, 0, 0, 0, 0, 1, 1),
		(drawing, 7497, 7497, 0, 0, 0, 0, 1, 1),
		(drawing, 7496, 7496, 0, 0, 0, 0, 1, 1),
		(drawing, 7495, 7495, 0, 0, 0, 0, 1, 1),
		(drawing, 7494, 7494, 0, 0, 0, 0, 1, 1),
		(drawing, 7493, 7493, 0, 0, 0, 0, 1, 1),
		(drawing, 7492, 7492, 0, 0, 0, 0, 1, 1),
		(drawing, 7491, 7491, 0, 0, 0, 0, 1, 1),
		(drawing, 7490, 7490, 0, 0, 0, 0, 1, 1),
		(drawing, 7489, 7489, 0, 0, 0, 0, 1, 1),
		(drawing, 7488, 7488, 0, 0, 0, 0, 1, 1),
		(drawing, 7487, 7487, 0, 0, 0, 0, 1, 1),
		(drawing, 7486, 7486, 0, 0, 0, 0, 1, 1),
		(drawing, 7485, 7485, 0, 0, 0, 0, 1, 1),
		(drawing, 7484, 7484, 0, 0, 0, 0, 1, 1),
		(drawing, 7483, 7483, 0, 0, 0, 0, 1, 1),
		(drawing, 7482, 7482, 0, 0, 0, 0, 1, 1),
		(drawing, 7481, 7481, 0, 0, 0, 0, 1, 1),
		(drawing, 7480, 7480, 0, 0, 0, 0, 1, 1),
		(drawing, 7479, 7479, 0, 0, 0, 0, 1, 1),
		(drawing, 7478, 7478, 0, 0, 0, 0, 1, 1),
		(drawing, 7477, 7477, 0, 0, 0, 0, 1, 1),
		(drawing, 7476, 7476, 0, 0, 0, 0, 1, 1),
		(drawing, 7475, 7475, 0, 0, 0, 0, 1, 1),
		(drawing, 7474, 7474, 0, 0, 0, 0, 1, 1),
		(drawing, 7473, 7473, 0, 0, 0, 0, 1, 1),
		(drawing, 7472, 7472, 0, 0, 0, 0, 1, 1),
		(drawing, 7471, 7471, 0, 0, 0, 0, 1, 1),
		(drawing, 7470, 7470, 0, 0, 0, 0, 1, 1),
		(drawing, 7469, 7469, 0, 0, 0, 0, 1, 1),
		(drawing, 7468, 7468, 0, 0, 0, 0, 1, 1),
		(drawing, 7467, 7467, 0, 0, 0, 0, 1, 1),
		(drawing, 7466, 7466, 0, 0, 0, 0, 1, 1),
		(drawing, 7465, 7465, 0, 0, 0, 0, 1, 1),
		(drawing, 7464, 7464, 0, 0, 0, 0, 1, 1),
		(drawing, 7463, 7463, 0, 0, 0, 0, 1, 1),
		(drawing, 7462, 7462, 0, 0, 0, 0, 1, 1),
		(drawing, 7461, 7461, 0, 0, 0, 0, 1, 1),
		(drawing, 7460, 7460, 0, 0, 0, 0, 1, 1),
		(drawing, 7459, 7459, 0, 0, 0, 0, 1, 1),
		(drawing, 7458, 7458, 0, 0, 0, 0, 1, 1),
		(drawing, 7457, 7457, 0, 0, 0, 0, 1, 1),
		(drawing, 7456, 7456, 0, 0, 0, 0, 1, 1),
		(drawing, 7455, 7455, 0, 0, 0, 0, 1, 1),
		(drawing, 7454, 7454, 0, 0, 0, 0, 1, 1),
		(drawing, 7453, 7453, 0, 0, 0, 0, 1, 1),
		(drawing, 7452, 7452, 0, 0, 0, 0, 1, 1),
		(drawing, 7451, 7451, 0, 0, 0, 0, 1, 1),
		(drawing, 7450, 7450, 0, 0, 0, 0, 1, 1),
		(drawing, 7449, 7449, 0, 0, 0, 0, 1, 1),
		(drawing, 7448, 7448, 0, 0, 0, 0, 1, 1),
		(drawing, 7447, 7447, 0, 0, 0, 0, 1, 1),
		(drawing, 7446, 7446, 0, 0, 0, 0, 1, 1),
		(drawing, 7445, 7445, 0, 0, 0, 0, 1, 1),
		(drawing, 7444, 7444, 0, 0, 0, 0, 1, 1),
		(drawing, 7443, 7443, 0, 0, 0, 0, 1, 1),
		(drawing, 7442, 7442, 0, 0, 0, 0, 1, 1),
		(drawing, 7441, 7441, 0, 0, 0, 0, 1, 1),
		(drawing, 7440, 7440, 0, 0, 0, 0, 1, 1),
		(drawing, 7439, 7439, 0, 0, 0, 0, 1, 1),
		(drawing, 7438, 7438, 0, 0, 0, 0, 1, 1),
		(drawing, 7437, 7437, 0, 0, 0, 0, 1, 1),
		(drawing, 7436, 7436, 0, 0, 0, 0, 1, 1),
		(drawing, 7435, 7435, 0, 0, 0, 0, 1, 1),
		(drawing, 7434, 7434, 0, 0, 0, 0, 1, 1),
		(drawing, 7433, 7433, 0, 0, 0, 0, 1, 1),
		(drawing, 7432, 7432, 0, 0, 0, 0, 1, 1),
		(drawing, 7431, 7431, 0, 0, 0, 0, 1, 1),
		(drawing, 7430, 7430, 0, 0, 0, 0, 1, 1),
		(drawing, 7429, 7429, 0, 0, 0, 0, 1, 1),
		(drawing, 7428, 7428, 0, 0, 0, 0, 1, 1),
		(drawing, 7427, 7427, 0, 0, 0, 0, 1, 1),
		(drawing, 7426, 7426, 0, 0, 0, 0, 1, 1),
		(drawing, 7425, 7425, 0, 0, 0, 0, 1, 1),
		(drawing, 7424, 7424, 0, 0, 0, 0, 1, 1),
		(drawing, 7423, 7423, 0, 0, 0, 0, 1, 1),
		(drawing, 7422, 7422, 0, 0, 0, 0, 1, 1),
		(drawing, 7421, 7421, 0, 0, 0, 0, 1, 1),
		(drawing, 7420, 7420, 0, 0, 0, 0, 1, 1),
		(drawing, 7419, 7419, 0, 0, 0, 0, 1, 1),
		(drawing, 7418, 7418, 0, 0, 0, 0, 1, 1),
		(drawing, 7417, 7417, 0, 0, 0, 0, 1, 1),
		(drawing, 7416, 7416, 0, 0, 0, 0, 1, 1),
		(drawing, 7415, 7415, 0, 0, 0, 0, 1, 1),
		(drawing, 7414, 7414, 0, 0, 0, 0, 1, 1),
		(drawing, 7413, 7413, 0, 0, 0, 0, 1, 1),
		(drawing, 7412, 7412, 0, 0, 0, 0, 1, 1),
		(drawing, 7411, 7411, 0, 0, 0, 0, 1, 1),
		(drawing, 7410, 7410, 0, 0, 0, 0, 1, 1),
		(drawing, 7409, 7409, 0, 0, 0, 0, 1, 1),
		(drawing, 7408, 7408, 0, 0, 0, 0, 1, 1),
		(drawing, 7407, 7407, 0, 0, 0, 0, 1, 1),
		(drawing, 7406, 7406, 0, 0, 0, 0, 1, 1),
		(drawing, 7405, 7405, 0, 0, 0, 0, 1, 1),
		(drawing, 7404, 7404, 0, 0, 0, 0, 1, 1),
		(drawing, 7403, 7403, 0, 0, 0, 0, 1, 1),
		(drawing, 7402, 7402, 0, 0, 0, 0, 1, 1),
		(drawing, 7401, 7401, 0, 0, 0, 0, 1, 1),
		(drawing, 7400, 7400, 0, 0, 0, 0, 1, 1),
		(drawing, 7399, 7399, 0, 0, 0, 0, 1, 1),
		(drawing, 7398, 7398, 0, 0, 0, 0, 1, 1),
		(drawing, 7397, 7397, 0, 0, 0, 0, 1, 1),
		(drawing, 7396, 7396, 0, 0, 0, 0, 1, 1),
		(drawing, 7395, 7395, 0, 0, 0, 0, 1, 1),
		(drawing, 7394, 7394, 0, 0, 0, 0, 1, 1),
		(drawing, 7393, 7393, 0, 0, 0, 0, 1, 1),
		(drawing, 7392, 7392, 0, 0, 0, 0, 1, 1),
		(drawing, 7391, 7391, 0, 0, 0, 0, 1, 1),
		(drawing, 7390, 7390, 0, 0, 0, 0, 1, 1),
		(drawing, 7389, 7389, 0, 0, 0, 0, 1, 1),
		(drawing, 7388, 7388, 0, 0, 0, 0, 1, 1),
		(drawing, 7387, 7387, 0, 0, 0, 0, 1, 1),
		(drawing, 7386, 7386, 0, 0, 0, 0, 1, 1),
		(drawing, 7385, 7385, 0, 0, 0, 0, 1, 1),
		(drawing, 7384, 7384, 0, 0, 0, 0, 1, 1),
		(drawing, 7383, 7383, 0, 0, 0, 0, 1, 1),
		(drawing, 7382, 7382, 0, 0, 0, 0, 1, 1),
		(drawing, 7381, 7381, 0, 0, 0, 0, 1, 1),
		(drawing, 7380, 7380, 0, 0, 0, 0, 1, 1),
		(drawing, 7379, 7379, 0, 0, 0, 0, 1, 1),
		(drawing, 7378, 7378, 0, 0, 0, 0, 1, 1),
		(drawing, 7377, 7377, 0, 0, 0, 0, 1, 1),
		(drawing, 7376, 7376, 0, 0, 0, 0, 1, 1),
		(drawing, 7375, 7375, 0, 0, 0, 0, 1, 1),
		(drawing, 7374, 7374, 0, 0, 0, 0, 1, 1),
		(drawing, 7373, 7373, 0, 0, 0, 0, 1, 1),
		(drawing, 7372, 7372, 0, 0, 0, 0, 1, 1),
		(drawing, 7371, 7371, 0, 0, 0, 0, 1, 1),
		(drawing, 7370, 7370, 0, 0, 0, 0, 1, 1),
		(drawing, 7369, 7369, 0, 0, 0, 0, 1, 1),
		(drawing, 7368, 7368, 0, 0, 0, 0, 1, 1),
		(drawing, 7367, 7367, 0, 0, 0, 0, 1, 1),
		(drawing, 7366, 7366, 0, 0, 0, 0, 1, 1),
		(drawing, 7365, 7365, 0, 0, 0, 0, 1, 1),
		(drawing, 7364, 7364, 0, 0, 0, 0, 1, 1),
		(drawing, 7363, 7363, 0, 0, 0, 0, 1, 1),
		(drawing, 7362, 7362, 0, 0, 0, 0, 1, 1),
		(drawing, 7361, 7361, 0, 0, 0, 0, 1, 1),
		(drawing, 7360, 7360, 0, 0, 0, 0, 1, 1),
		(drawing, 7359, 7359, 0, 0, 0, 0, 1, 1),
		(drawing, 7358, 7358, 0, 0, 0, 0, 1, 1),
		(drawing, 7357, 7357, 0, 0, 0, 0, 1, 1),
		(drawing, 7356, 7356, 0, 0, 0, 0, 1, 1),
		(drawing, 7355, 7355, 0, 0, 0, 0, 1, 1),
		(drawing, 7354, 7354, 0, 0, 0, 0, 1, 1),
		(drawing, 7353, 7353, 0, 0, 0, 0, 1, 1),
		(drawing, 7352, 7352, 0, 0, 0, 0, 1, 1),
		(drawing, 7351, 7351, 0, 0, 0, 0, 1, 1),
		(drawing, 7350, 7350, 0, 0, 0, 0, 1, 1),
		(drawing, 7349, 7349, 0, 0, 0, 0, 1, 1),
		(drawing, 7348, 7348, 0, 0, 0, 0, 1, 1),
		(drawing, 7347, 7347, 0, 0, 0, 0, 1, 1),
		(drawing, 7346, 7346, 0, 0, 0, 0, 1, 1),
		(drawing, 7345, 7345, 0, 0, 0, 0, 1, 1),
		(drawing, 7344, 7344, 0, 0, 0, 0, 1, 1),
		(drawing, 7343, 7343, 0, 0, 0, 0, 1, 1),
		(drawing, 7342, 7342, 0, 0, 0, 0, 1, 1),
		(drawing, 7341, 7341, 0, 0, 0, 0, 1, 1),
		(drawing, 7340, 7340, 0, 0, 0, 0, 1, 1),
		(drawing, 7339, 7339, 0, 0, 0, 0, 1, 1),
		(drawing, 7338, 7338, 0, 0, 0, 0, 1, 1),
		(drawing, 7337, 7337, 0, 0, 0, 0, 1, 1),
		(drawing, 7336, 7336, 0, 0, 0, 0, 1, 1),
		(drawing, 7335, 7335, 0, 0, 0, 0, 1, 1),
		(drawing, 7334, 7334, 0, 0, 0, 0, 1, 1),
		(drawing, 7333, 7333, 0, 0, 0, 0, 1, 1),
		(drawing, 7332, 7332, 0, 0, 0, 0, 1, 1),
		(drawing, 7331, 7331, 0, 0, 0, 0, 1, 1),
		(drawing, 7330, 7330, 0, 0, 0, 0, 1, 1),
		(drawing, 7329, 7329, 0, 0, 0, 0, 1, 1),
		(drawing, 7328, 7328, 0, 0, 0, 0, 1, 1),
		(drawing, 7327, 7327, 0, 0, 0, 0, 1, 1),
		(drawing, 7326, 7326, 0, 0, 0, 0, 1, 1),
		(drawing, 7325, 7325, 0, 0, 0, 0, 1, 1),
		(drawing, 7324, 7324, 0, 0, 0, 0, 1, 1),
		(drawing, 7323, 7323, 0, 0, 0, 0, 1, 1),
		(drawing, 7322, 7322, 0, 0, 0, 0, 1, 1),
		(drawing, 7321, 7321, 0, 0, 0, 0, 1, 1),
		(drawing, 7320, 7320, 0, 0, 0, 0, 1, 1),
		(drawing, 7319, 7319, 0, 0, 0, 0, 1, 1),
		(drawing, 7318, 7318, 0, 0, 0, 0, 1, 1),
		(drawing, 7317, 7317, 0, 0, 0, 0, 1, 1),
		(drawing, 7316, 7316, 0, 0, 0, 0, 1, 1),
		(drawing, 7315, 7315, 0, 0, 0, 0, 1, 1),
		(drawing, 7314, 7314, 0, 0, 0, 0, 1, 1),
		(drawing, 7313, 7313, 0, 0, 0, 0, 1, 1),
		(drawing, 7312, 7312, 0, 0, 0, 0, 1, 1),
		(drawing, 7311, 7311, 0, 0, 0, 0, 1, 1),
		(drawing, 7310, 7310, 0, 0, 0, 0, 1, 1),
		(drawing, 7309, 7309, 0, 0, 0, 0, 1, 1),
		(drawing, 7308, 7308, 0, 0, 0, 0, 1, 1),
		(drawing, 7307, 7307, 0, 0, 0, 0, 1, 1),
		(drawing, 7306, 7306, 0, 0, 0, 0, 1, 1),
		(drawing, 7305, 7305, 0, 0, 0, 0, 1, 1),
		(drawing, 7304, 7304, 0, 0, 0, 0, 1, 1),
		(drawing, 7303, 7303, 0, 0, 0, 0, 1, 1),
		(drawing, 7302, 7302, 0, 0, 0, 0, 1, 1),
		(drawing, 7301, 7301, 0, 0, 0, 0, 1, 1),
		(drawing, 7300, 7300, 0, 0, 0, 0, 1, 1),
		(drawing, 7299, 7299, 0, 0, 0, 0, 1, 1),
		(drawing, 7298, 7298, 0, 0, 0, 0, 1, 1),
		(drawing, 7297, 7297, 0, 0, 0, 0, 1, 1),
		(drawing, 7296, 7296, 0, 0, 0, 0, 1, 1),
		(drawing, 7295, 7295, 0, 0, 0, 0, 1, 1),
		(drawing, 7294, 7294, 0, 0, 0, 0, 1, 1),
		(drawing, 7293, 7293, 0, 0, 0, 0, 1, 1),
		(drawing, 7292, 7292, 0, 0, 0, 0, 1, 1),
		(drawing, 7291, 7291, 0, 0, 0, 0, 1, 1),
		(drawing, 7290, 7290, 0, 0, 0, 0, 1, 1),
		(drawing, 7289, 7289, 0, 0, 0, 0, 1, 1),
		(drawing, 7288, 7288, 0, 0, 0, 0, 1, 1),
		(drawing, 7287, 7287, 0, 0, 0, 0, 1, 1),
		(drawing, 7286, 7286, 0, 0, 0, 0, 1, 1),
		(drawing, 7285, 7285, 0, 0, 0, 0, 1, 1),
		(drawing, 7284, 7284, 0, 0, 0, 0, 1, 1),
		(drawing, 7283, 7283, 0, 0, 0, 0, 1, 1),
		(drawing, 7282, 7282, 0, 0, 0, 0, 1, 1),
		(drawing, 7281, 7281, 0, 0, 0, 0, 1, 1),
		(drawing, 7280, 7280, 0, 0, 0, 0, 1, 1),
		(drawing, 7279, 7279, 0, 0, 0, 0, 1, 1),
		(drawing, 7278, 7278, 0, 0, 0, 0, 1, 1),
		(drawing, 7277, 7277, 0, 0, 0, 0, 1, 1),
		(drawing, 7276, 7276, 0, 0, 0, 0, 1, 1),
		(drawing, 7275, 7275, 0, 0, 0, 0, 1, 1),
		(drawing, 7274, 7274, 0, 0, 0, 0, 1, 1),
		(drawing, 7273, 7273, 0, 0, 0, 0, 1, 1),
		(drawing, 7272, 7272, 0, 0, 0, 0, 1, 1),
		(drawing, 7271, 7271, 0, 0, 0, 0, 1, 1),
		(drawing, 7270, 7270, 0, 0, 0, 0, 1, 1),
		(drawing, 7269, 7269, 0, 0, 0, 0, 1, 1),
		(drawing, 7268, 7268, 0, 0, 0, 0, 1, 1),
		(drawing, 7267, 7267, 0, 0, 0, 0, 1, 1),
		(drawing, 7266, 7266, 0, 0, 0, 0, 1, 1),
		(drawing, 7265, 7265, 0, 0, 0, 0, 1, 1),
		(drawing, 7264, 7264, 0, 0, 0, 0, 1, 1),
		(drawing, 7263, 7263, 0, 0, 0, 0, 1, 1),
		(drawing, 7262, 7262, 0, 0, 0, 0, 1, 1),
		(drawing, 7261, 7261, 0, 0, 0, 0, 1, 1),
		(drawing, 7260, 7260, 0, 0, 0, 0, 1, 1),
		(drawing, 7259, 7259, 0, 0, 0, 0, 1, 1),
		(drawing, 7258, 7258, 0, 0, 0, 0, 1, 1),
		(drawing, 7257, 7257, 0, 0, 0, 0, 1, 1),
		(drawing, 7256, 7256, 0, 0, 0, 0, 1, 1),
		(drawing, 7255, 7255, 0, 0, 0, 0, 1, 1),
		(drawing, 7254, 7254, 0, 0, 0, 0, 1, 1),
		(drawing, 7253, 7253, 0, 0, 0, 0, 1, 1),
		(drawing, 7252, 7252, 0, 0, 0, 0, 1, 1),
		(drawing, 7251, 7251, 0, 0, 0, 0, 1, 1),
		(drawing, 7250, 7250, 0, 0, 0, 0, 1, 1),
		(drawing, 7249, 7249, 0, 0, 0, 0, 1, 1),
		(drawing, 7248, 7248, 0, 0, 0, 0, 1, 1),
		(drawing, 7247, 7247, 0, 0, 0, 0, 1, 1),
		(drawing, 7246, 7246, 0, 0, 0, 0, 1, 1),
		(drawing, 7245, 7245, 0, 0, 0, 0, 1, 1),
		(drawing, 7244, 7244, 0, 0, 0, 0, 1, 1),
		(drawing, 7243, 7243, 0, 0, 0, 0, 1, 1),
		(drawing, 7242, 7242, 0, 0, 0, 0, 1, 1),
		(drawing, 7241, 7241, 0, 0, 0, 0, 1, 1),
		(drawing, 7240, 7240, 0, 0, 0, 0, 1, 1),
		(drawing, 7239, 7239, 0, 0, 0, 0, 1, 1),
		(drawing, 7238, 7238, 0, 0, 0, 0, 1, 1),
		(drawing, 7237, 7237, 0, 0, 0, 0, 1, 1),
		(drawing, 7236, 7236, 0, 0, 0, 0, 1, 1),
		(drawing, 7235, 7235, 0, 0, 0, 0, 1, 1),
		(drawing, 7234, 7234, 0, 0, 0, 0, 1, 1),
		(drawing, 7233, 7233, 0, 0, 0, 0, 1, 1),
		(drawing, 7232, 7232, 0, 0, 0, 0, 1, 1),
		(drawing, 7231, 7231, 0, 0, 0, 0, 1, 1),
		(drawing, 7230, 7230, 0, 0, 0, 0, 1, 1),
		(drawing, 7229, 7229, 0, 0, 0, 0, 1, 1),
		(drawing, 7228, 7228, 0, 0, 0, 0, 1, 1),
		(drawing, 7227, 7227, 0, 0, 0, 0, 1, 1),
		(drawing, 7226, 7226, 0, 0, 0, 0, 1, 1),
		(drawing, 7225, 7225, 0, 0, 0, 0, 1, 1),
		(drawing, 7224, 7224, 0, 0, 0, 0, 1, 1),
		(drawing, 7223, 7223, 0, 0, 0, 0, 1, 1),
		(drawing, 7222, 7222, 0, 0, 0, 0, 1, 1),
		(drawing, 7221, 7221, 0, 0, 0, 0, 1, 1),
		(drawing, 7220, 7220, 0, 0, 0, 0, 1, 1),
		(drawing, 7219, 7219, 0, 0, 0, 0, 1, 1),
		(drawing, 7218, 7218, 0, 0, 0, 0, 1, 1),
		(drawing, 7217, 7217, 0, 0, 0, 0, 1, 1),
		(drawing, 7216, 7216, 0, 0, 0, 0, 1, 1),
		(drawing, 7215, 7215, 0, 0, 0, 0, 1, 1),
		(drawing, 7214, 7214, 0, 0, 0, 0, 1, 1),
		(drawing, 7213, 7213, 0, 0, 0, 0, 1, 1),
		(drawing, 7212, 7212, 0, 0, 0, 0, 1, 1),
		(drawing, 7211, 7211, 0, 0, 0, 0, 1, 1),
		(drawing, 7210, 7210, 0, 0, 0, 0, 1, 1),
		(drawing, 7209, 7209, 0, 0, 0, 0, 1, 1),
		(drawing, 7208, 7208, 0, 0, 0, 0, 1, 1),
		(drawing, 7207, 7207, 0, 0, 0, 0, 1, 1),
		(drawing, 7206, 7206, 0, 0, 0, 0, 1, 1),
		(drawing, 7205, 7205, 0, 0, 0, 0, 1, 1),
		(drawing, 7204, 7204, 0, 0, 0, 0, 1, 1),
		(drawing, 7203, 7203, 0, 0, 0, 0, 1, 1),
		(drawing, 7202, 7202, 0, 0, 0, 0, 1, 1),
		(drawing, 7201, 7201, 0, 0, 0, 0, 1, 1),
		(drawing, 7200, 7200, 0, 0, 0, 0, 1, 1),
		(drawing, 7199, 7199, 0, 0, 0, 0, 1, 1),
		(drawing, 7198, 7198, 0, 0, 0, 0, 1, 1),
		(drawing, 7197, 7197, 0, 0, 0, 0, 1, 1),
		(drawing, 7196, 7196, 0, 0, 0, 0, 1, 1),
		(drawing, 7195, 7195, 0, 0, 0, 0, 1, 1),
		(drawing, 7194, 7194, 0, 0, 0, 0, 1, 1),
		(drawing, 7193, 7193, 0, 0, 0, 0, 1, 1),
		(drawing, 7192, 7192, 0, 0, 0, 0, 1, 1),
		(drawing, 7191, 7191, 0, 0, 0, 0, 1, 1),
		(drawing, 7190, 7190, 0, 0, 0, 0, 1, 1),
		(drawing, 7189, 7189, 0, 0, 0, 0, 1, 1),
		(drawing, 7188, 7188, 0, 0, 0, 0, 1, 1),
		(drawing, 7187, 7187, 0, 0, 0, 0, 1, 1),
		(drawing, 7186, 7186, 0, 0, 0, 0, 1, 1),
		(drawing, 7185, 7185, 0, 0, 0, 0, 1, 1),
		(drawing, 7184, 7184, 0, 0, 0, 0, 1, 1),
		(drawing, 7183, 7183, 0, 0, 0, 0, 1, 1),
		(drawing, 7182, 7182, 0, 0, 0, 0, 1, 1),
		(drawing, 7181, 7181, 0, 0, 0, 0, 1, 1),
		(drawing, 7180, 7180, 0, 0, 0, 0, 1, 1),
		(drawing, 7179, 7179, 0, 0, 0, 0, 1, 1),
		(drawing, 7178, 7178, 0, 0, 0, 0, 1, 1),
		(drawing, 7177, 7177, 0, 0, 0, 0, 1, 1),
		(drawing, 7176, 7176, 0, 0, 0, 0, 1, 1),
		(drawing, 7175, 7175, 0, 0, 0, 0, 1, 1),
		(drawing, 7174, 7174, 0, 0, 0, 0, 1, 1),
		(drawing, 7173, 7173, 0, 0, 0, 0, 1, 1),
		(drawing, 7172, 7172, 0, 0, 0, 0, 1, 1),
		(drawing, 7171, 7171, 0, 0, 0, 0, 1, 1),
		(drawing, 7170, 7170, 0, 0, 0, 0, 1, 1),
		(drawing, 7169, 7169, 0, 0, 0, 0, 1, 1),
		(drawing, 7168, 7168, 0, 0, 0, 0, 1, 1),
		(drawing, 7167, 7167, 0, 0, 0, 0, 1, 1),
		(drawing, 7166, 7166, 0, 0, 0, 0, 1, 1),
		(drawing, 7165, 7165, 0, 0, 0, 0, 1, 1),
		(drawing, 7164, 7164, 0, 0, 0, 0, 1, 1),
		(drawing, 7163, 7163, 0, 0, 0, 0, 1, 1),
		(drawing, 7162, 7162, 0, 0, 0, 0, 1, 1),
		(drawing, 7161, 7161, 0, 0, 0, 0, 1, 1),
		(drawing, 7160, 7160, 0, 0, 0, 0, 1, 1),
		(drawing, 7159, 7159, 0, 0, 0, 0, 1, 1),
		(drawing, 7158, 7158, 0, 0, 0, 0, 1, 1),
		(drawing, 7157, 7157, 0, 0, 0, 0, 1, 1),
		(drawing, 7156, 7156, 0, 0, 0, 0, 1, 1),
		(drawing, 7155, 7155, 0, 0, 0, 0, 1, 1),
		(drawing, 7154, 7154, 0, 0, 0, 0, 1, 1),
		(drawing, 7153, 7153, 0, 0, 0, 0, 1, 1),
		(drawing, 7152, 7152, 0, 0, 0, 0, 1, 1),
		(drawing, 7151, 7151, 0, 0, 0, 0, 1, 1),
		(drawing, 7150, 7150, 0, 0, 0, 0, 1, 1),
		(drawing, 7149, 7149, 0, 0, 0, 0, 1, 1),
		(drawing, 7148, 7148, 0, 0, 0, 0, 1, 1),
		(drawing, 7147, 7147, 0, 0, 0, 0, 1, 1),
		(drawing, 7146, 7146, 0, 0, 0, 0, 1, 1),
		(drawing, 7145, 7145, 0, 0, 0, 0, 1, 1),
		(drawing, 7144, 7144, 0, 0, 0, 0, 1, 1),
		(drawing, 7143, 7143, 0, 0, 0, 0, 1, 1),
		(drawing, 7142, 7142, 0, 0, 0, 0, 1, 1),
		(drawing, 7141, 7141, 0, 0, 0, 0, 1, 1),
		(drawing, 7140, 7140, 0, 0, 0, 0, 1, 1),
		(drawing, 7139, 7139, 0, 0, 0, 0, 1, 1),
		(drawing, 7138, 7138, 0, 0, 0, 0, 1, 1),
		(drawing, 7137, 7137, 0, 0, 0, 0, 1, 1),
		(drawing, 7136, 7136, 0, 0, 0, 0, 1, 1),
		(drawing, 7135, 7135, 0, 0, 0, 0, 1, 1),
		(drawing, 7134, 7134, 0, 0, 0, 0, 1, 1),
		(drawing, 7133, 7133, 0, 0, 0, 0, 1, 1),
		(drawing, 7132, 7132, 0, 0, 0, 0, 1, 1),
		(drawing, 7131, 7131, 0, 0, 0, 0, 1, 1),
		(drawing, 7130, 7130, 0, 0, 0, 0, 1, 1),
		(drawing, 7129, 7129, 0, 0, 0, 0, 1, 1),
		(drawing, 7128, 7128, 0, 0, 0, 0, 1, 1),
		(drawing, 7127, 7127, 0, 0, 0, 0, 1, 1),
		(drawing, 7126, 7126, 0, 0, 0, 0, 1, 1),
		(drawing, 7125, 7125, 0, 0, 0, 0, 1, 1),
		(drawing, 7124, 7124, 0, 0, 0, 0, 1, 1),
		(drawing, 7123, 7123, 0, 0, 0, 0, 1, 1),
		(drawing, 7122, 7122, 0, 0, 0, 0, 1, 1),
		(drawing, 7121, 7121, 0, 0, 0, 0, 1, 1),
		(drawing, 7120, 7120, 0, 0, 0, 0, 1, 1),
		(drawing, 7119, 7119, 0, 0, 0, 0, 1, 1),
		(drawing, 7118, 7118, 0, 0, 0, 0, 1, 1),
		(drawing, 7117, 7117, 0, 0, 0, 0, 1, 1),
		(drawing, 7116, 7116, 0, 0, 0, 0, 1, 1),
		(drawing, 7115, 7115, 0, 0, 0, 0, 1, 1),
		(drawing, 7114, 7114, 0, 0, 0, 0, 1, 1),
		(drawing, 7113, 7113, 0, 0, 0, 0, 1, 1),
		(drawing, 7112, 7112, 0, 0, 0, 0, 1, 1),
		(drawing, 7111, 7111, 0, 0, 0, 0, 1, 1),
		(drawing, 7110, 7110, 0, 0, 0, 0, 1, 1),
		(drawing, 7109, 7109, 0, 0, 0, 0, 1, 1),
		(drawing, 7108, 7108, 0, 0, 0, 0, 1, 1),
		(drawing, 7107, 7107, 0, 0, 0, 0, 1, 1),
		(drawing, 7106, 7106, 0, 0, 0, 0, 1, 1),
		(drawing, 7105, 7105, 0, 0, 0, 0, 1, 1),
		(drawing, 7104, 7104, 0, 0, 0, 0, 1, 1),
		(drawing, 7103, 7103, 0, 0, 0, 0, 1, 1),
		(drawing, 7102, 7102, 0, 0, 0, 0, 1, 1),
		(drawing, 7101, 7101, 0, 0, 0, 0, 1, 1),
		(drawing, 7100, 7100, 0, 0, 0, 0, 1, 1),
		(drawing, 7099, 7099, 0, 0, 0, 0, 1, 1),
		(drawing, 7098, 7098, 0, 0, 0, 0, 1, 1),
		(drawing, 7097, 7097, 0, 0, 0, 0, 1, 1),
		(drawing, 7096, 7096, 0, 0, 0, 0, 1, 1),
		(drawing, 7095, 7095, 0, 0, 0, 0, 1, 1),
		(drawing, 7094, 7094, 0, 0, 0, 0, 1, 1),
		(drawing, 7093, 7093, 0, 0, 0, 0, 1, 1),
		(drawing, 7092, 7092, 0, 0, 0, 0, 1, 1),
		(drawing, 7091, 7091, 0, 0, 0, 0, 1, 1),
		(drawing, 7090, 7090, 0, 0, 0, 0, 1, 1),
		(drawing, 7089, 7089, 0, 0, 0, 0, 1, 1),
		(drawing, 7088, 7088, 0, 0, 0, 0, 1, 1),
		(drawing, 7087, 7087, 0, 0, 0, 0, 1, 1),
		(drawing, 7086, 7086, 0, 0, 0, 0, 1, 1),
		(drawing, 7085, 7085, 0, 0, 0, 0, 1, 1),
		(drawing, 7084, 7084, 0, 0, 0, 0, 1, 1),
		(drawing, 7083, 7083, 0, 0, 0, 0, 1, 1),
		(drawing, 7082, 7082, 0, 0, 0, 0, 1, 1),
		(drawing, 7081, 7081, 0, 0, 0, 0, 1, 1),
		(drawing, 7080, 7080, 0, 0, 0, 0, 1, 1),
		(drawing, 7079, 7079, 0, 0, 0, 0, 1, 1),
		(drawing, 7078, 7078, 0, 0, 0, 0, 1, 1),
		(drawing, 7077, 7077, 0, 0, 0, 0, 1, 1),
		(drawing, 7076, 7076, 0, 0, 0, 0, 1, 1),
		(drawing, 7075, 7075, 0, 0, 0, 0, 1, 1),
		(drawing, 7074, 7074, 0, 0, 0, 0, 1, 1),
		(drawing, 7073, 7073, 0, 0, 0, 0, 1, 1),
		(drawing, 7072, 7072, 0, 0, 0, 0, 1, 1),
		(drawing, 7071, 7071, 0, 0, 0, 0, 1, 1),
		(drawing, 7070, 7070, 0, 0, 0, 0, 1, 1),
		(drawing, 7069, 7069, 0, 0, 0, 0, 1, 1),
		(drawing, 7068, 7068, 0, 0, 0, 0, 1, 1),
		(drawing, 7067, 7067, 0, 0, 0, 0, 1, 1),
		(drawing, 7066, 7066, 0, 0, 0, 0, 1, 1),
		(drawing, 7065, 7065, 0, 0, 0, 0, 1, 1),
		(drawing, 7064, 7064, 0, 0, 0, 0, 1, 1),
		(drawing, 7063, 7063, 0, 0, 0, 0, 1, 1),
		(drawing, 7062, 7062, 0, 0, 0, 0, 1, 1),
		(drawing, 7061, 7061, 0, 0, 0, 0, 1, 1),
		(drawing, 7060, 7060, 0, 0, 0, 0, 1, 1),
		(drawing, 7059, 7059, 0, 0, 0, 0, 1, 1),
		(drawing, 7058, 7058, 0, 0, 0, 0, 1, 1),
		(drawing, 7057, 7057, 0, 0, 0, 0, 1, 1),
		(drawing, 7056, 7056, 0, 0, 0, 0, 1, 1),
		(drawing, 7055, 7055, 0, 0, 0, 0, 1, 1),
		(drawing, 7054, 7054, 0, 0, 0, 0, 1, 1),
		(drawing, 7053, 7053, 0, 0, 0, 0, 1, 1),
		(drawing, 7052, 7052, 0, 0, 0, 0, 1, 1),
		(drawing, 7051, 7051, 0, 0, 0, 0, 1, 1),
		(drawing, 7050, 7050, 0, 0, 0, 0, 1, 1),
		(drawing, 7049, 7049, 0, 0, 0, 0, 1, 1),
		(drawing, 7048, 7048, 0, 0, 0, 0, 1, 1),
		(drawing, 7047, 7047, 0, 0, 0, 0, 1, 1),
		(drawing, 7046, 7046, 0, 0, 0, 0, 1, 1),
		(drawing, 7045, 7045, 0, 0, 0, 0, 1, 1),
		(drawing, 7044, 7044, 0, 0, 0, 0, 1, 1),
		(drawing, 7043, 7043, 0, 0, 0, 0, 1, 1),
		(drawing, 7042, 7042, 0, 0, 0, 0, 1, 1),
		(drawing, 7041, 7041, 0, 0, 0, 0, 1, 1),
		(drawing, 7040, 7040, 0, 0, 0, 0, 1, 1),
		(drawing, 7039, 7039, 0, 0, 0, 0, 1, 1),
		(drawing, 7038, 7038, 0, 0, 0, 0, 1, 1),
		(drawing, 7037, 7037, 0, 0, 0, 0, 1, 1),
		(drawing, 7036, 7036, 0, 0, 0, 0, 1, 1),
		(drawing, 7035, 7035, 0, 0, 0, 0, 1, 1),
		(drawing, 7034, 7034, 0, 0, 0, 0, 1, 1),
		(drawing, 7033, 7033, 0, 0, 0, 0, 1, 1),
		(drawing, 7032, 7032, 0, 0, 0, 0, 1, 1),
		(drawing, 7031, 7031, 0, 0, 0, 0, 1, 1),
		(drawing, 7030, 7030, 0, 0, 0, 0, 1, 1),
		(drawing, 7029, 7029, 0, 0, 0, 0, 1, 1),
		(drawing, 7028, 7028, 0, 0, 0, 0, 1, 1),
		(drawing, 7027, 7027, 0, 0, 0, 0, 1, 1),
		(drawing, 7026, 7026, 0, 0, 0, 0, 1, 1),
		(drawing, 7025, 7025, 0, 0, 0, 0, 1, 1),
		(drawing, 7024, 7024, 0, 0, 0, 0, 1, 1),
		(drawing, 7023, 7023, 0, 0, 0, 0, 1, 1),
		(drawing, 7022, 7022, 0, 0, 0, 0, 1, 1),
		(drawing, 7021, 7021, 0, 0, 0, 0, 1, 1),
		(drawing, 7020, 7020, 0, 0, 0, 0, 1, 1),
		(drawing, 7019, 7019, 0, 0, 0, 0, 1, 1),
		(drawing, 7018, 7018, 0, 0, 0, 0, 1, 1),
		(drawing, 7017, 7017, 0, 0, 0, 0, 1, 1),
		(drawing, 7016, 7016, 0, 0, 0, 0, 1, 1),
		(drawing, 7015, 7015, 0, 0, 0, 0, 1, 1),
		(drawing, 7014, 7014, 0, 0, 0, 0, 1, 1),
		(drawing, 7013, 7013, 0, 0, 0, 0, 1, 1),
		(drawing, 7012, 7012, 0, 0, 0, 0, 1, 1),
		(drawing, 7011, 7011, 0, 0, 0, 0, 1, 1),
		(drawing, 7010, 7010, 0, 0, 0, 0, 1, 1),
		(drawing, 7009, 7009, 0, 0, 0, 0, 1, 1),
		(drawing, 7008, 7008, 0, 0, 0, 0, 1, 1),
		(drawing, 7007, 7007, 0, 0, 0, 0, 1, 1),
		(drawing, 7006, 7006, 0, 0, 0, 0, 1, 1),
		(drawing, 7005, 7005, 0, 0, 0, 0, 1, 1),
		(drawing, 7004, 7004, 0, 0, 0, 0, 1, 1),
		(drawing, 7003, 7003, 0, 0, 0, 0, 1, 1),
		(drawing, 7002, 7002, 0, 0, 0, 0, 1, 1),
		(drawing, 7001, 7001, 0, 0, 0, 0, 1, 1),
		(drawing, 7000, 7000, 0, 0, 0, 0, 1, 1),
		(drawing, 6999, 6999, 0, 0, 0, 0, 1, 1),
		(drawing, 6998, 6998, 0, 0, 0, 0, 1, 1),
		(drawing, 6997, 6997, 0, 0, 0, 0, 1, 1),
		(drawing, 6996, 6996, 0, 0, 0, 0, 1, 1),
		(drawing, 6995, 6995, 0, 0, 0, 0, 1, 1),
		(drawing, 6994, 6994, 0, 0, 0, 0, 1, 1),
		(drawing, 6993, 6993, 0, 0, 0, 0, 1, 1),
		(drawing, 6992, 6992, 0, 0, 0, 0, 1, 1),
		(drawing, 6991, 6991, 0, 0, 0, 0, 1, 1),
		(drawing, 6990, 6990, 0, 0, 0, 0, 1, 1),
		(drawing, 6989, 6989, 0, 0, 0, 0, 1, 1),
		(drawing, 6988, 6988, 0, 0, 0, 0, 1, 1),
		(drawing, 6987, 6987, 0, 0, 0, 0, 1, 1),
		(drawing, 6986, 6986, 0, 0, 0, 0, 1, 1),
		(drawing, 6985, 6985, 0, 0, 0, 0, 1, 1),
		(drawing, 6984, 6984, 0, 0, 0, 0, 1, 1),
		(drawing, 6983, 6983, 0, 0, 0, 0, 1, 1),
		(drawing, 6982, 6982, 0, 0, 0, 0, 1, 1),
		(drawing, 6981, 6981, 0, 0, 0, 0, 1, 1),
		(drawing, 6980, 6980, 0, 0, 0, 0, 1, 1),
		(drawing, 6979, 6979, 0, 0, 0, 0, 1, 1),
		(drawing, 6978, 6978, 0, 0, 0, 0, 1, 1),
		(drawing, 6977, 6977, 0, 0, 0, 0, 1, 1),
		(drawing, 6976, 6976, 0, 0, 0, 0, 1, 1),
		(drawing, 6975, 6975, 0, 0, 0, 0, 1, 1),
		(drawing, 6974, 6974, 0, 0, 0, 0, 1, 1),
		(drawing, 6973, 6973, 0, 0, 0, 0, 1, 1),
		(drawing, 6972, 6972, 0, 0, 0, 0, 1, 1),
		(drawing, 6971, 6971, 0, 0, 0, 0, 1, 1),
		(drawing, 6970, 6970, 0, 0, 0, 0, 1, 1),
		(drawing, 6969, 6969, 0, 0, 0, 0, 1, 1),
		(drawing, 6968, 6968, 0, 0, 0, 0, 1, 1),
		(drawing, 6967, 6967, 0, 0, 0, 0, 1, 1),
		(drawing, 6966, 6966, 0, 0, 0, 0, 1, 1),
		(drawing, 6965, 6965, 0, 0, 0, 0, 1, 1),
		(drawing, 6964, 6964, 0, 0, 0, 0, 1, 1),
		(drawing, 6963, 6963, 0, 0, 0, 0, 1, 1),
		(drawing, 6962, 6962, 0, 0, 0, 0, 1, 1),
		(drawing, 6961, 6961, 0, 0, 0, 0, 1, 1),
		(drawing, 6960, 6960, 0, 0, 0, 0, 1, 1),
		(drawing, 6959, 6959, 0, 0, 0, 0, 1, 1),
		(drawing, 6958, 6958, 0, 0, 0, 0, 1, 1),
		(drawing, 6957, 6957, 0, 0, 0, 0, 1, 1),
		(drawing, 6956, 6956, 0, 0, 0, 0, 1, 1),
		(drawing, 6955, 6955, 0, 0, 0, 0, 1, 1),
		(drawing, 6954, 6954, 0, 0, 0, 0, 1, 1),
		(drawing, 6953, 6953, 0, 0, 0, 0, 1, 1),
		(drawing, 6952, 6952, 0, 0, 0, 0, 1, 1),
		(drawing, 6951, 6951, 0, 0, 0, 0, 1, 1),
		(drawing, 6950, 6950, 0, 0, 0, 0, 1, 1),
		(drawing, 6949, 6949, 0, 0, 0, 0, 1, 1),
		(drawing, 6948, 6948, 0, 0, 0, 0, 1, 1),
		(drawing, 6947, 6947, 0, 0, 0, 0, 1, 1),
		(drawing, 6946, 6946, 0, 0, 0, 0, 1, 1),
		(drawing, 6945, 6945, 0, 0, 0, 0, 1, 1),
		(drawing, 6944, 6944, 0, 0, 0, 0, 1, 1),
		(drawing, 6943, 6943, 0, 0, 0, 0, 1, 1),
		(drawing, 6942, 6942, 0, 0, 0, 0, 1, 1),
		(drawing, 6941, 6941, 0, 0, 0, 0, 1, 1),
		(drawing, 6940, 6940, 0, 0, 0, 0, 1, 1),
		(drawing, 6939, 6939, 0, 0, 0, 0, 1, 1),
		(drawing, 6938, 6938, 0, 0, 0, 0, 1, 1),
		(drawing, 6937, 6937, 0, 0, 0, 0, 1, 1),
		(drawing, 6936, 6936, 0, 0, 0, 0, 1, 1),
		(drawing, 6935, 6935, 0, 0, 0, 0, 1, 1),
		(drawing, 6934, 6934, 0, 0, 0, 0, 1, 1),
		(drawing, 6933, 6933, 0, 0, 0, 0, 1, 1),
		(drawing, 6932, 6932, 0, 0, 0, 0, 1, 1),
		(drawing, 6931, 6931, 0, 0, 0, 0, 1, 1),
		(drawing, 6930, 6930, 0, 0, 0, 0, 1, 1),
		(drawing, 6929, 6929, 0, 0, 0, 0, 1, 1),
		(drawing, 6928, 6928, 0, 0, 0, 0, 1, 1),
		(drawing, 6927, 6927, 0, 0, 0, 0, 1, 1),
		(drawing, 6926, 6926, 0, 0, 0, 0, 1, 1),
		(drawing, 6925, 6925, 0, 0, 0, 0, 1, 1),
		(drawing, 6924, 6924, 0, 0, 0, 0, 1, 1),
		(drawing, 6923, 6923, 0, 0, 0, 0, 1, 1),
		(drawing, 6922, 6922, 0, 0, 0, 0, 1, 1),
		(drawing, 6921, 6921, 0, 0, 0, 0, 1, 1),
		(drawing, 6920, 6920, 0, 0, 0, 0, 1, 1),
		(drawing, 6919, 6919, 0, 0, 0, 0, 1, 1),
		(drawing, 6918, 6918, 0, 0, 0, 0, 1, 1),
		(drawing, 6917, 6917, 0, 0, 0, 0, 1, 1),
		(drawing, 6916, 6916, 0, 0, 0, 0, 1, 1),
		(drawing, 6915, 6915, 0, 0, 0, 0, 1, 1),
		(drawing, 6914, 6914, 0, 0, 0, 0, 1, 1),
		(drawing, 6913, 6913, 0, 0, 0, 0, 1, 1),
		(drawing, 6912, 6912, 0, 0, 0, 0, 1, 1),
		(drawing, 6911, 6911, 0, 0, 0, 0, 1, 1),
		(drawing, 6910, 6910, 0, 0, 0, 0, 1, 1),
		(drawing, 6909, 6909, 0, 0, 0, 0, 1, 1),
		(drawing, 6908, 6908, 0, 0, 0, 0, 1, 1),
		(drawing, 6907, 6907, 0, 0, 0, 0, 1, 1),
		(drawing, 6906, 6906, 0, 0, 0, 0, 1, 1),
		(drawing, 6905, 6905, 0, 0, 0, 0, 1, 1),
		(drawing, 6904, 6904, 0, 0, 0, 0, 1, 1),
		(drawing, 6903, 6903, 0, 0, 0, 0, 1, 1),
		(drawing, 6902, 6902, 0, 0, 0, 0, 1, 1),
		(drawing, 6901, 6901, 0, 0, 0, 0, 1, 1),
		(drawing, 6900, 6900, 0, 0, 0, 0, 1, 1),
		(drawing, 6899, 6899, 0, 0, 0, 0, 1, 1),
		(drawing, 6898, 6898, 0, 0, 0, 0, 1, 1),
		(drawing, 6897, 6897, 0, 0, 0, 0, 1, 1),
		(drawing, 6896, 6896, 0, 0, 0, 0, 1, 1),
		(drawing, 6895, 6895, 0, 0, 0, 0, 1, 1),
		(drawing, 6894, 6894, 0, 0, 0, 0, 1, 1),
		(drawing, 6893, 6893, 0, 0, 0, 0, 1, 1),
		(drawing, 6892, 6892, 0, 0, 0, 0, 1, 1),
		(drawing, 6891, 6891, 0, 0, 0, 0, 1, 1),
		(drawing, 6890, 6890, 0, 0, 0, 0, 1, 1),
		(drawing, 6889, 6889, 0, 0, 0, 0, 1, 1),
		(drawing, 6888, 6888, 0, 0, 0, 0, 1, 1),
		(drawing, 6887, 6887, 0, 0, 0, 0, 1, 1),
		(drawing, 6886, 6886, 0, 0, 0, 0, 1, 1),
		(drawing, 6885, 6885, 0, 0, 0, 0, 1, 1),
		(drawing, 6884, 6884, 0, 0, 0, 0, 1, 1),
		(drawing, 6883, 6883, 0, 0, 0, 0, 1, 1),
		(drawing, 6882, 6882, 0, 0, 0, 0, 1, 1),
		(drawing, 6881, 6881, 0, 0, 0, 0, 1, 1),
		(drawing, 6880, 6880, 0, 0, 0, 0, 1, 1),
		(drawing, 6879, 6879, 0, 0, 0, 0, 1, 1),
		(drawing, 6878, 6878, 0, 0, 0, 0, 1, 1),
		(drawing, 6877, 6877, 0, 0, 0, 0, 1, 1),
		(drawing, 6876, 6876, 0, 0, 0, 0, 1, 1),
		(drawing, 6875, 6875, 0, 0, 0, 0, 1, 1),
		(drawing, 6874, 6874, 0, 0, 0, 0, 1, 1),
		(drawing, 6873, 6873, 0, 0, 0, 0, 1, 1),
		(drawing, 6872, 6872, 0, 0, 0, 0, 1, 1),
		(drawing, 6871, 6871, 0, 0, 0, 0, 1, 1),
		(drawing, 6870, 6870, 0, 0, 0, 0, 1, 1),
		(drawing, 6869, 6869, 0, 0, 0, 0, 1, 1),
		(drawing, 6868, 6868, 0, 0, 0, 0, 1, 1),
		(drawing, 6867, 6867, 0, 0, 0, 0, 1, 1),
		(drawing, 6866, 6866, 0, 0, 0, 0, 1, 1),
		(drawing, 6865, 6865, 0, 0, 0, 0, 1, 1),
		(drawing, 6864, 6864, 0, 0, 0, 0, 1, 1),
		(drawing, 6863, 6863, 0, 0, 0, 0, 1, 1),
		(drawing, 6862, 6862, 0, 0, 0, 0, 1, 1),
		(drawing, 6861, 6861, 0, 0, 0, 0, 1, 1),
		(drawing, 6860, 6860, 0, 0, 0, 0, 1, 1),
		(drawing, 6859, 6859, 0, 0, 0, 0, 1, 1),
		(drawing, 6858, 6858, 0, 0, 0, 0, 1, 1),
		(drawing, 6857, 6857, 0, 0, 0, 0, 1, 1),
		(drawing, 6856, 6856, 0, 0, 0, 0, 1, 1),
		(drawing, 6855, 6855, 0, 0, 0, 0, 1, 1),
		(drawing, 6854, 6854, 0, 0, 0, 0, 1, 1),
		(drawing, 6853, 6853, 0, 0, 0, 0, 1, 1),
		(drawing, 6852, 6852, 0, 0, 0, 0, 1, 1),
		(drawing, 6851, 6851, 0, 0, 0, 0, 1, 1),
		(drawing, 6850, 6850, 0, 0, 0, 0, 1, 1),
		(drawing, 6849, 6849, 0, 0, 0, 0, 1, 1),
		(drawing, 6848, 6848, 0, 0, 0, 0, 1, 1),
		(drawing, 6847, 6847, 0, 0, 0, 0, 1, 1),
		(drawing, 6846, 6846, 0, 0, 0, 0, 1, 1),
		(drawing, 6845, 6845, 0, 0, 0, 0, 1, 1),
		(drawing, 6844, 6844, 0, 0, 0, 0, 1, 1),
		(drawing, 6843, 6843, 0, 0, 0, 0, 1, 1),
		(drawing, 6842, 6842, 0, 0, 0, 0, 1, 1),
		(drawing, 6841, 6841, 0, 0, 0, 0, 1, 1),
		(drawing, 6840, 6840, 0, 0, 0, 0, 1, 1),
		(drawing, 6839, 6839, 0, 0, 0, 0, 1, 1),
		(drawing, 6838, 6838, 0, 0, 0, 0, 1, 1),
		(drawing, 6837, 6837, 0, 0, 0, 0, 1, 1),
		(drawing, 6836, 6836, 0, 0, 0, 0, 1, 1),
		(drawing, 6835, 6835, 0, 0, 0, 0, 1, 1),
		(drawing, 6834, 6834, 0, 0, 0, 0, 1, 1),
		(drawing, 6833, 6833, 0, 0, 0, 0, 1, 1),
		(drawing, 6832, 6832, 0, 0, 0, 0, 1, 1),
		(drawing, 6831, 6831, 0, 0, 0, 0, 1, 1),
		(drawing, 6830, 6830, 0, 0, 0, 0, 1, 1),
		(drawing, 6829, 6829, 0, 0, 0, 0, 1, 1),
		(drawing, 6828, 6828, 0, 0, 0, 0, 1, 1),
		(drawing, 6827, 6827, 0, 0, 0, 0, 1, 1),
		(drawing, 6826, 6826, 0, 0, 0, 0, 1, 1),
		(drawing, 6825, 6825, 0, 0, 0, 0, 1, 1),
		(drawing, 6824, 6824, 0, 0, 0, 0, 1, 1),
		(drawing, 6823, 6823, 0, 0, 0, 0, 1, 1),
		(drawing, 6822, 6822, 0, 0, 0, 0, 1, 1),
		(drawing, 6821, 6821, 0, 0, 0, 0, 1, 1),
		(drawing, 6820, 6820, 0, 0, 0, 0, 1, 1),
		(drawing, 6819, 6819, 0, 0, 0, 0, 1, 1),
		(drawing, 6818, 6818, 0, 0, 0, 0, 1, 1),
		(drawing, 6817, 6817, 0, 0, 0, 0, 1, 1),
		(drawing, 6816, 6816, 0, 0, 0, 0, 1, 1),
		(drawing, 6815, 6815, 0, 0, 0, 0, 1, 1),
		(drawing, 6814, 6814, 0, 0, 0, 0, 1, 1),
		(drawing, 6813, 6813, 0, 0, 0, 0, 1, 1),
		(drawing, 6812, 6812, 0, 0, 0, 0, 1, 1),
		(drawing, 6811, 6811, 0, 0, 0, 0, 1, 1),
		(drawing, 6810, 6810, 0, 0, 0, 0, 1, 1),
		(drawing, 6809, 6809, 0, 0, 0, 0, 1, 1),
		(drawing, 6808, 6808, 0, 0, 0, 0, 1, 1),
		(drawing, 6807, 6807, 0, 0, 0, 0, 1, 1),
		(drawing, 6806, 6806, 0, 0, 0, 0, 1, 1),
		(drawing, 6805, 6805, 0, 0, 0, 0, 1, 1),
		(drawing, 6804, 6804, 0, 0, 0, 0, 1, 1),
		(drawing, 6803, 6803, 0, 0, 0, 0, 1, 1),
		(drawing, 6802, 6802, 0, 0, 0, 0, 1, 1),
		(drawing, 6801, 6801, 0, 0, 0, 0, 1, 1),
		(drawing, 6800, 6800, 0, 0, 0, 0, 1, 1),
		(drawing, 6799, 6799, 0, 0, 0, 0, 1, 1),
		(drawing, 6798, 6798, 0, 0, 0, 0, 1, 1),
		(drawing, 6797, 6797, 0, 0, 0, 0, 1, 1),
		(drawing, 6796, 6796, 0, 0, 0, 0, 1, 1),
		(drawing, 6795, 6795, 0, 0, 0, 0, 1, 1),
		(drawing, 6794, 6794, 0, 0, 0, 0, 1, 1),
		(drawing, 6793, 6793, 0, 0, 0, 0, 1, 1),
		(drawing, 6792, 6792, 0, 0, 0, 0, 1, 1),
		(drawing, 6791, 6791, 0, 0, 0, 0, 1, 1),
		(drawing, 6790, 6790, 0, 0, 0, 0, 1, 1),
		(drawing, 6789, 6789, 0, 0, 0, 0, 1, 1),
		(drawing, 6788, 6788, 0, 0, 0, 0, 1, 1),
		(drawing, 6787, 6787, 0, 0, 0, 0, 1, 1),
		(drawing, 6786, 6786, 0, 0, 0, 0, 1, 1),
		(drawing, 6785, 6785, 0, 0, 0, 0, 1, 1),
		(drawing, 6784, 6784, 0, 0, 0, 0, 1, 1),
		(drawing, 6783, 6783, 0, 0, 0, 0, 1, 1),
		(drawing, 6782, 6782, 0, 0, 0, 0, 1, 1),
		(drawing, 6781, 6781, 0, 0, 0, 0, 1, 1),
		(drawing, 6780, 6780, 0, 0, 0, 0, 1, 1),
		(drawing, 6779, 6779, 0, 0, 0, 0, 1, 1),
		(drawing, 6778, 6778, 0, 0, 0, 0, 1, 1),
		(drawing, 6777, 6777, 0, 0, 0, 0, 1, 1),
		(drawing, 6776, 6776, 0, 0, 0, 0, 1, 1),
		(drawing, 6775, 6775, 0, 0, 0, 0, 1, 1),
		(drawing, 6774, 6774, 0, 0, 0, 0, 1, 1),
		(drawing, 6773, 6773, 0, 0, 0, 0, 1, 1),
		(drawing, 6772, 6772, 0, 0, 0, 0, 1, 1),
		(drawing, 6771, 6771, 0, 0, 0, 0, 1, 1),
		(drawing, 6770, 6770, 0, 0, 0, 0, 1, 1),
		(drawing, 6769, 6769, 0, 0, 0, 0, 1, 1),
		(drawing, 6768, 6768, 0, 0, 0, 0, 1, 1),
		(drawing, 6767, 6767, 0, 0, 0, 0, 1, 1),
		(drawing, 6766, 6766, 0, 0, 0, 0, 1, 1),
		(drawing, 6765, 6765, 0, 0, 0, 0, 1, 1),
		(drawing, 6764, 6764, 0, 0, 0, 0, 1, 1),
		(drawing, 6763, 6763, 0, 0, 0, 0, 1, 1),
		(drawing, 6762, 6762, 0, 0, 0, 0, 1, 1),
		(drawing, 6761, 6761, 0, 0, 0, 0, 1, 1),
		(drawing, 6760, 6760, 0, 0, 0, 0, 1, 1),
		(drawing, 6759, 6759, 0, 0, 0, 0, 1, 1),
		(drawing, 6758, 6758, 0, 0, 0, 0, 1, 1),
		(drawing, 6757, 6757, 0, 0, 0, 0, 1, 1),
		(drawing, 6756, 6756, 0, 0, 0, 0, 1, 1),
		(drawing, 6755, 6755, 0, 0, 0, 0, 1, 1),
		(drawing, 6754, 6754, 0, 0, 0, 0, 1, 1),
		(drawing, 6753, 6753, 0, 0, 0, 0, 1, 1),
		(drawing, 6752, 6752, 0, 0, 0, 0, 1, 1),
		(drawing, 6751, 6751, 0, 0, 0, 0, 1, 1),
		(drawing, 6750, 6750, 0, 0, 0, 0, 1, 1),
		(drawing, 6749, 6749, 0, 0, 0, 0, 1, 1),
		(drawing, 6748, 6748, 0, 0, 0, 0, 1, 1),
		(drawing, 6747, 6747, 0, 0, 0, 0, 1, 1),
		(drawing, 6746, 6746, 0, 0, 0, 0, 1, 1),
		(drawing, 6745, 6745, 0, 0, 0, 0, 1, 1),
		(drawing, 6744, 6744, 0, 0, 0, 0, 1, 1),
		(drawing, 6743, 6743, 0, 0, 0, 0, 1, 1),
		(drawing, 6742, 6742, 0, 0, 0, 0, 1, 1),
		(drawing, 6741, 6741, 0, 0, 0, 0, 1, 1),
		(drawing, 6740, 6740, 0, 0, 0, 0, 1, 1),
		(drawing, 6739, 6739, 0, 0, 0, 0, 1, 1),
		(drawing, 6738, 6738, 0, 0, 0, 0, 1, 1),
		(drawing, 6737, 6737, 0, 0, 0, 0, 1, 1),
		(drawing, 6736, 6736, 0, 0, 0, 0, 1, 1),
		(drawing, 6735, 6735, 0, 0, 0, 0, 1, 1),
		(drawing, 6734, 6734, 0, 0, 0, 0, 1, 1),
		(drawing, 6733, 6733, 0, 0, 0, 0, 1, 1),
		(drawing, 6732, 6732, 0, 0, 0, 0, 1, 1),
		(drawing, 6731, 6731, 0, 0, 0, 0, 1, 1),
		(drawing, 6730, 6730, 0, 0, 0, 0, 1, 1),
		(drawing, 6729, 6729, 0, 0, 0, 0, 1, 1),
		(drawing, 6728, 6728, 0, 0, 0, 0, 1, 1),
		(drawing, 6727, 6727, 0, 0, 0, 0, 1, 1),
		(drawing, 6726, 6726, 0, 0, 0, 0, 1, 1),
		(drawing, 6725, 6725, 0, 0, 0, 0, 1, 1),
		(drawing, 6724, 6724, 0, 0, 0, 0, 1, 1),
		(drawing, 6723, 6723, 0, 0, 0, 0, 1, 1),
		(drawing, 6722, 6722, 0, 0, 0, 0, 1, 1),
		(drawing, 6721, 6721, 0, 0, 0, 0, 1, 1),
		(drawing, 6720, 6720, 0, 0, 0, 0, 1, 1),
		(drawing, 6719, 6719, 0, 0, 0, 0, 1, 1),
		(drawing, 6718, 6718, 0, 0, 0, 0, 1, 1),
		(drawing, 6717, 6717, 0, 0, 0, 0, 1, 1),
		(drawing, 6716, 6716, 0, 0, 0, 0, 1, 1),
		(drawing, 6715, 6715, 0, 0, 0, 0, 1, 1),
		(drawing, 6714, 6714, 0, 0, 0, 0, 1, 1),
		(drawing, 6713, 6713, 0, 0, 0, 0, 1, 1),
		(drawing, 6712, 6712, 0, 0, 0, 0, 1, 1),
		(drawing, 6711, 6711, 0, 0, 0, 0, 1, 1),
		(drawing, 6710, 6710, 0, 0, 0, 0, 1, 1),
		(drawing, 6709, 6709, 0, 0, 0, 0, 1, 1),
		(drawing, 6708, 6708, 0, 0, 0, 0, 1, 1),
		(drawing, 6707, 6707, 0, 0, 0, 0, 1, 1),
		(drawing, 6706, 6706, 0, 0, 0, 0, 1, 1),
		(drawing, 6705, 6705, 0, 0, 0, 0, 1, 1),
		(drawing, 6704, 6704, 0, 0, 0, 0, 1, 1),
		(drawing, 6703, 6703, 0, 0, 0, 0, 1, 1),
		(drawing, 6702, 6702, 0, 0, 0, 0, 1, 1),
		(drawing, 6701, 6701, 0, 0, 0, 0, 1, 1),
		(drawing, 6700, 6700, 0, 0, 0, 0, 1, 1),
		(drawing, 6699, 6699, 0, 0, 0, 0, 1, 1),
		(drawing, 6698, 6698, 0, 0, 0, 0, 1, 1),
		(drawing, 6697, 6697, 0, 0, 0, 0, 1, 1),
		(drawing, 6696, 6696, 0, 0, 0, 0, 1, 1),
		(drawing, 6695, 6695, 0, 0, 0, 0, 1, 1),
		(drawing, 6694, 6694, 0, 0, 0, 0, 1, 1),
		(drawing, 6693, 6693, 0, 0, 0, 0, 1, 1),
		(drawing, 6692, 6692, 0, 0, 0, 0, 1, 1),
		(drawing, 6691, 6691, 0, 0, 0, 0, 1, 1),
		(drawing, 6690, 6690, 0, 0, 0, 0, 1, 1),
		(drawing, 6689, 6689, 0, 0, 0, 0, 1, 1),
		(drawing, 6688, 6688, 0, 0, 0, 0, 1, 1),
		(drawing, 6687, 6687, 0, 0, 0, 0, 1, 1),
		(drawing, 6686, 6686, 0, 0, 0, 0, 1, 1),
		(drawing, 6685, 6685, 0, 0, 0, 0, 1, 1),
		(drawing, 6684, 6684, 0, 0, 0, 0, 1, 1),
		(drawing, 6683, 6683, 0, 0, 0, 0, 1, 1),
		(drawing, 6682, 6682, 0, 0, 0, 0, 1, 1),
		(drawing, 6681, 6681, 0, 0, 0, 0, 1, 1),
		(drawing, 6680, 6680, 0, 0, 0, 0, 1, 1),
		(drawing, 6679, 6679, 0, 0, 0, 0, 1, 1),
		(drawing, 6678, 6678, 0, 0, 0, 0, 1, 1),
		(drawing, 6677, 6677, 0, 0, 0, 0, 1, 1),
		(drawing, 6676, 6676, 0, 0, 0, 0, 1, 1),
		(drawing, 6675, 6675, 0, 0, 0, 0, 1, 1),
		(drawing, 6674, 6674, 0, 0, 0, 0, 1, 1),
		(drawing, 6673, 6673, 0, 0, 0, 0, 1, 1),
		(drawing, 6672, 6672, 0, 0, 0, 0, 1, 1),
		(drawing, 6671, 6671, 0, 0, 0, 0, 1, 1),
		(drawing, 6670, 6670, 0, 0, 0, 0, 1, 1),
		(drawing, 6669, 6669, 0, 0, 0, 0, 1, 1),
		(drawing, 6668, 6668, 0, 0, 0, 0, 1, 1),
		(drawing, 6667, 6667, 0, 0, 0, 0, 1, 1),
		(drawing, 6666, 6666, 0, 0, 0, 0, 1, 1),
		(drawing, 6665, 6665, 0, 0, 0, 0, 1, 1),
		(drawing, 6664, 6664, 0, 0, 0, 0, 1, 1),
		(drawing, 6663, 6663, 0, 0, 0, 0, 1, 1),
		(drawing, 6662, 6662, 0, 0, 0, 0, 1, 1),
		(drawing, 6661, 6661, 0, 0, 0, 0, 1, 1),
		(drawing, 6660, 6660, 0, 0, 0, 0, 1, 1),
		(drawing, 6659, 6659, 0, 0, 0, 0, 1, 1),
		(drawing, 6658, 6658, 0, 0, 0, 0, 1, 1),
		(drawing, 6657, 6657, 0, 0, 0, 0, 1, 1),
		(drawing, 6656, 6656, 0, 0, 0, 0, 1, 1),
		(drawing, 6655, 6655, 0, 0, 0, 0, 1, 1),
		(drawing, 6654, 6654, 0, 0, 0, 0, 1, 1),
		(drawing, 6653, 6653, 0, 0, 0, 0, 1, 1),
		(drawing, 6652, 6652, 0, 0, 0, 0, 1, 1),
		(drawing, 6651, 6651, 0, 0, 0, 0, 1, 1),
		(drawing, 6650, 6650, 0, 0, 0, 0, 1, 1),
		(drawing, 6649, 6649, 0, 0, 0, 0, 1, 1),
		(drawing, 6648, 6648, 0, 0, 0, 0, 1, 1),
		(drawing, 6647, 6647, 0, 0, 0, 0, 1, 1),
		(drawing, 6646, 6646, 0, 0, 0, 0, 1, 1),
		(drawing, 6645, 6645, 0, 0, 0, 0, 1, 1),
		(drawing, 6644, 6644, 0, 0, 0, 0, 1, 1),
		(drawing, 6643, 6643, 0, 0, 0, 0, 1, 1),
		(drawing, 6642, 6642, 0, 0, 0, 0, 1, 1),
		(drawing, 6641, 6641, 0, 0, 0, 0, 1, 1),
		(drawing, 6640, 6640, 0, 0, 0, 0, 1, 1),
		(drawing, 6639, 6639, 0, 0, 0, 0, 1, 1),
		(drawing, 6638, 6638, 0, 0, 0, 0, 1, 1),
		(drawing, 6637, 6637, 0, 0, 0, 0, 1, 1),
		(drawing, 6636, 6636, 0, 0, 0, 0, 1, 1),
		(drawing, 6635, 6635, 0, 0, 0, 0, 1, 1),
		(drawing, 6634, 6634, 0, 0, 0, 0, 1, 1),
		(drawing, 6633, 6633, 0, 0, 0, 0, 1, 1),
		(drawing, 6632, 6632, 0, 0, 0, 0, 1, 1),
		(drawing, 6631, 6631, 0, 0, 0, 0, 1, 1),
		(drawing, 6630, 6630, 0, 0, 0, 0, 1, 1),
		(drawing, 6629, 6629, 0, 0, 0, 0, 1, 1),
		(drawing, 6628, 6628, 0, 0, 0, 0, 1, 1),
		(drawing, 6627, 6627, 0, 0, 0, 0, 1, 1),
		(drawing, 6626, 6626, 0, 0, 0, 0, 1, 1),
		(drawing, 6625, 6625, 0, 0, 0, 0, 1, 1),
		(drawing, 6624, 6624, 0, 0, 0, 0, 1, 1),
		(drawing, 6623, 6623, 0, 0, 0, 0, 1, 1),
		(drawing, 6622, 6622, 0, 0, 0, 0, 1, 1),
		(drawing, 6621, 6621, 0, 0, 0, 0, 1, 1),
		(drawing, 6620, 6620, 0, 0, 0, 0, 1, 1),
		(drawing, 6619, 6619, 0, 0, 0, 0, 1, 1),
		(drawing, 6618, 6618, 0, 0, 0, 0, 1, 1),
		(drawing, 6617, 6617, 0, 0, 0, 0, 1, 1),
		(drawing, 6616, 6616, 0, 0, 0, 0, 1, 1),
		(drawing, 6615, 6615, 0, 0, 0, 0, 1, 1),
		(drawing, 6614, 6614, 0, 0, 0, 0, 1, 1),
		(drawing, 6613, 6613, 0, 0, 0, 0, 1, 1),
		(drawing, 6612, 6612, 0, 0, 0, 0, 1, 1),
		(drawing, 6611, 6611, 0, 0, 0, 0, 1, 1),
		(drawing, 6610, 6610, 0, 0, 0, 0, 1, 1),
		(drawing, 6609, 6609, 0, 0, 0, 0, 1, 1),
		(drawing, 6608, 6608, 0, 0, 0, 0, 1, 1),
		(drawing, 6607, 6607, 0, 0, 0, 0, 1, 1),
		(drawing, 6606, 6606, 0, 0, 0, 0, 1, 1),
		(drawing, 6605, 6605, 0, 0, 0, 0, 1, 1),
		(drawing, 6604, 6604, 0, 0, 0, 0, 1, 1),
		(drawing, 6603, 6603, 0, 0, 0, 0, 1, 1),
		(drawing, 6602, 6602, 0, 0, 0, 0, 1, 1),
		(drawing, 6601, 6601, 0, 0, 0, 0, 1, 1),
		(drawing, 6600, 6600, 0, 0, 0, 0, 1, 1),
		(drawing, 6599, 6599, 0, 0, 0, 0, 1, 1),
		(drawing, 6598, 6598, 0, 0, 0, 0, 1, 1),
		(drawing, 6597, 6597, 0, 0, 0, 0, 1, 1),
		(drawing, 6596, 6596, 0, 0, 0, 0, 1, 1),
		(drawing, 6595, 6595, 0, 0, 0, 0, 1, 1),
		(drawing, 6594, 6594, 0, 0, 0, 0, 1, 1),
		(drawing, 6593, 6593, 0, 0, 0, 0, 1, 1),
		(drawing, 6592, 6592, 0, 0, 0, 0, 1, 1),
		(drawing, 6591, 6591, 0, 0, 0, 0, 1, 1),
		(drawing, 6590, 6590, 0, 0, 0, 0, 1, 1),
		(drawing, 6589, 6589, 0, 0, 0, 0, 1, 1),
		(drawing, 6588, 6588, 0, 0, 0, 0, 1, 1),
		(drawing, 6587, 6587, 0, 0, 0, 0, 1, 1),
		(drawing, 6586, 6586, 0, 0, 0, 0, 1, 1),
		(drawing, 6585, 6585, 0, 0, 0, 0, 1, 1),
		(drawing, 6584, 6584, 0, 0, 0, 0, 1, 1),
		(drawing, 6583, 6583, 0, 0, 0, 0, 1, 1),
		(drawing, 6582, 6582, 0, 0, 0, 0, 1, 1),
		(drawing, 6581, 6581, 0, 0, 0, 0, 1, 1),
		(drawing, 6580, 6580, 0, 0, 0, 0, 1, 1),
		(drawing, 6579, 6579, 0, 0, 0, 0, 1, 1),
		(drawing, 6578, 6578, 0, 0, 0, 0, 1, 1),
		(drawing, 6577, 6577, 0, 0, 0, 0, 1, 1),
		(drawing, 6576, 6576, 0, 0, 0, 0, 1, 1),
		(drawing, 6575, 6575, 0, 0, 0, 0, 1, 1),
		(drawing, 6574, 6574, 0, 0, 0, 0, 1, 1),
		(drawing, 6573, 6573, 0, 0, 0, 0, 1, 1),
		(drawing, 6572, 6572, 0, 0, 0, 0, 1, 1),
		(drawing, 6571, 6571, 0, 0, 0, 0, 1, 1),
		(drawing, 6570, 6570, 0, 0, 0, 0, 1, 1),
		(drawing, 6569, 6569, 0, 0, 0, 0, 1, 1),
		(drawing, 6568, 6568, 0, 0, 0, 0, 1, 1),
		(drawing, 6567, 6567, 0, 0, 0, 0, 1, 1),
		(drawing, 6566, 6566, 0, 0, 0, 0, 1, 1),
		(drawing, 6565, 6565, 0, 0, 0, 0, 1, 1),
		(drawing, 6564, 6564, 0, 0, 0, 0, 1, 1),
		(drawing, 6563, 6563, 0, 0, 0, 0, 1, 1),
		(drawing, 6562, 6562, 0, 0, 0, 0, 1, 1),
		(drawing, 6561, 6561, 0, 0, 0, 0, 1, 1),
		(drawing, 6560, 6560, 0, 0, 0, 0, 1, 1),
		(drawing, 6559, 6559, 0, 0, 0, 0, 1, 1),
		(drawing, 6558, 6558, 0, 0, 0, 0, 1, 1),
		(drawing, 6557, 6557, 0, 0, 0, 0, 1, 1),
		(drawing, 6556, 6556, 0, 0, 0, 0, 1, 1),
		(drawing, 6555, 6555, 0, 0, 0, 0, 1, 1),
		(drawing, 6554, 6554, 0, 0, 0, 0, 1, 1),
		(drawing, 6553, 6553, 0, 0, 0, 0, 1, 1),
		(drawing, 6552, 6552, 0, 0, 0, 0, 1, 1),
		(drawing, 6551, 6551, 0, 0, 0, 0, 1, 1),
		(drawing, 6550, 6550, 0, 0, 0, 0, 1, 1),
		(drawing, 6549, 6549, 0, 0, 0, 0, 1, 1),
		(drawing, 6548, 6548, 0, 0, 0, 0, 1, 1),
		(drawing, 6547, 6547, 0, 0, 0, 0, 1, 1),
		(drawing, 6546, 6546, 0, 0, 0, 0, 1, 1),
		(drawing, 6545, 6545, 0, 0, 0, 0, 1, 1),
		(drawing, 6544, 6544, 0, 0, 0, 0, 1, 1),
		(drawing, 6543, 6543, 0, 0, 0, 0, 1, 1),
		(drawing, 6542, 6542, 0, 0, 0, 0, 1, 1),
		(drawing, 6541, 6541, 0, 0, 0, 0, 1, 1),
		(drawing, 6540, 6540, 0, 0, 0, 0, 1, 1),
		(drawing, 6539, 6539, 0, 0, 0, 0, 1, 1),
		(drawing, 6538, 6538, 0, 0, 0, 0, 1, 1),
		(drawing, 6537, 6537, 0, 0, 0, 0, 1, 1),
		(drawing, 6536, 6536, 0, 0, 0, 0, 1, 1),
		(drawing, 6535, 6535, 0, 0, 0, 0, 1, 1),
		(drawing, 6534, 6534, 0, 0, 0, 0, 1, 1),
		(drawing, 6533, 6533, 0, 0, 0, 0, 1, 1),
		(drawing, 6532, 6532, 0, 0, 0, 0, 1, 1),
		(drawing, 6531, 6531, 0, 0, 0, 0, 1, 1),
		(drawing, 6530, 6530, 0, 0, 0, 0, 1, 1),
		(drawing, 6529, 6529, 0, 0, 0, 0, 1, 1),
		(drawing, 6528, 6528, 0, 0, 0, 0, 1, 1),
		(drawing, 6527, 6527, 0, 0, 0, 0, 1, 1),
		(drawing, 6526, 6526, 0, 0, 0, 0, 1, 1),
		(drawing, 6525, 6525, 0, 0, 0, 0, 1, 1),
		(drawing, 6524, 6524, 0, 0, 0, 0, 1, 1),
		(drawing, 6523, 6523, 0, 0, 0, 0, 1, 1),
		(drawing, 6522, 6522, 0, 0, 0, 0, 1, 1),
		(drawing, 6521, 6521, 0, 0, 0, 0, 1, 1),
		(drawing, 6520, 6520, 0, 0, 0, 0, 1, 1),
		(drawing, 6519, 6519, 0, 0, 0, 0, 1, 1),
		(drawing, 6518, 6518, 0, 0, 0, 0, 1, 1),
		(drawing, 6517, 6517, 0, 0, 0, 0, 1, 1),
		(drawing, 6516, 6516, 0, 0, 0, 0, 1, 1),
		(drawing, 6515, 6515, 0, 0, 0, 0, 1, 1),
		(drawing, 6514, 6514, 0, 0, 0, 0, 1, 1),
		(drawing, 6513, 6513, 0, 0, 0, 0, 1, 1),
		(drawing, 6512, 6512, 0, 0, 0, 0, 1, 1),
		(drawing, 6511, 6511, 0, 0, 0, 0, 1, 1),
		(drawing, 6510, 6510, 0, 0, 0, 0, 1, 1),
		(drawing, 6509, 6509, 0, 0, 0, 0, 1, 1),
		(drawing, 6508, 6508, 0, 0, 0, 0, 1, 1),
		(drawing, 6507, 6507, 0, 0, 0, 0, 1, 1),
		(drawing, 6506, 6506, 0, 0, 0, 0, 1, 1),
		(drawing, 6505, 6505, 0, 0, 0, 0, 1, 1),
		(drawing, 6504, 6504, 0, 0, 0, 0, 1, 1),
		(drawing, 6503, 6503, 0, 0, 0, 0, 1, 1),
		(drawing, 6502, 6502, 0, 0, 0, 0, 1, 1),
		(drawing, 6501, 6501, 0, 0, 0, 0, 1, 1),
		(drawing, 6500, 6500, 0, 0, 0, 0, 1, 1),
		(drawing, 6499, 6499, 0, 0, 0, 0, 1, 1),
		(drawing, 6498, 6498, 0, 0, 0, 0, 1, 1),
		(drawing, 6497, 6497, 0, 0, 0, 0, 1, 1),
		(drawing, 6496, 6496, 0, 0, 0, 0, 1, 1),
		(drawing, 6495, 6495, 0, 0, 0, 0, 1, 1),
		(drawing, 6494, 6494, 0, 0, 0, 0, 1, 1),
		(drawing, 6493, 6493, 0, 0, 0, 0, 1, 1),
		(drawing, 6492, 6492, 0, 0, 0, 0, 1, 1),
		(drawing, 6491, 6491, 0, 0, 0, 0, 1, 1),
		(drawing, 6490, 6490, 0, 0, 0, 0, 1, 1),
		(drawing, 6489, 6489, 0, 0, 0, 0, 1, 1),
		(drawing, 6488, 6488, 0, 0, 0, 0, 1, 1),
		(drawing, 6487, 6487, 0, 0, 0, 0, 1, 1),
		(drawing, 6486, 6486, 0, 0, 0, 0, 1, 1),
		(drawing, 6485, 6485, 0, 0, 0, 0, 1, 1),
		(drawing, 6484, 6484, 0, 0, 0, 0, 1, 1),
		(drawing, 6483, 6483, 0, 0, 0, 0, 1, 1),
		(drawing, 6482, 6482, 0, 0, 0, 0, 1, 1),
		(drawing, 6481, 6481, 0, 0, 0, 0, 1, 1),
		(drawing, 6480, 6480, 0, 0, 0, 0, 1, 1),
		(drawing, 6479, 6479, 0, 0, 0, 0, 1, 1),
		(drawing, 6478, 6478, 0, 0, 0, 0, 1, 1),
		(drawing, 6477, 6477, 0, 0, 0, 0, 1, 1),
		(drawing, 6476, 6476, 0, 0, 0, 0, 1, 1),
		(drawing, 6475, 6475, 0, 0, 0, 0, 1, 1),
		(drawing, 6474, 6474, 0, 0, 0, 0, 1, 1),
		(drawing, 6473, 6473, 0, 0, 0, 0, 1, 1),
		(drawing, 6472, 6472, 0, 0, 0, 0, 1, 1),
		(drawing, 6471, 6471, 0, 0, 0, 0, 1, 1),
		(drawing, 6470, 6470, 0, 0, 0, 0, 1, 1),
		(drawing, 6469, 6469, 0, 0, 0, 0, 1, 1),
		(drawing, 6468, 6468, 0, 0, 0, 0, 1, 1),
		(drawing, 6467, 6467, 0, 0, 0, 0, 1, 1),
		(drawing, 6466, 6466, 0, 0, 0, 0, 1, 1),
		(drawing, 6465, 6465, 0, 0, 0, 0, 1, 1),
		(drawing, 6464, 6464, 0, 0, 0, 0, 1, 1),
		(drawing, 6463, 6463, 0, 0, 0, 0, 1, 1),
		(drawing, 6462, 6462, 0, 0, 0, 0, 1, 1),
		(drawing, 6461, 6461, 0, 0, 0, 0, 1, 1),
		(drawing, 6460, 6460, 0, 0, 0, 0, 1, 1),
		(drawing, 6459, 6459, 0, 0, 0, 0, 1, 1),
		(drawing, 6458, 6458, 0, 0, 0, 0, 1, 1),
		(drawing, 6457, 6457, 0, 0, 0, 0, 1, 1),
		(drawing, 6456, 6456, 0, 0, 0, 0, 1, 1),
		(drawing, 6455, 6455, 0, 0, 0, 0, 1, 1),
		(drawing, 6454, 6454, 0, 0, 0, 0, 1, 1),
		(drawing, 6453, 6453, 0, 0, 0, 0, 1, 1),
		(drawing, 6452, 6452, 0, 0, 0, 0, 1, 1),
		(drawing, 6451, 6451, 0, 0, 0, 0, 1, 1),
		(drawing, 6450, 6450, 0, 0, 0, 0, 1, 1),
		(drawing, 6449, 6449, 0, 0, 0, 0, 1, 1),
		(drawing, 6448, 6448, 0, 0, 0, 0, 1, 1),
		(drawing, 6447, 6447, 0, 0, 0, 0, 1, 1),
		(drawing, 6446, 6446, 0, 0, 0, 0, 1, 1),
		(drawing, 6445, 6445, 0, 0, 0, 0, 1, 1),
		(drawing, 6444, 6444, 0, 0, 0, 0, 1, 1),
		(drawing, 6443, 6443, 0, 0, 0, 0, 1, 1),
		(drawing, 6442, 6442, 0, 0, 0, 0, 1, 1),
		(drawing, 6441, 6441, 0, 0, 0, 0, 1, 1),
		(drawing, 6440, 6440, 0, 0, 0, 0, 1, 1),
		(drawing, 6439, 6439, 0, 0, 0, 0, 1, 1),
		(drawing, 6438, 6438, 0, 0, 0, 0, 1, 1),
		(drawing, 6437, 6437, 0, 0, 0, 0, 1, 1),
		(drawing, 6436, 6436, 0, 0, 0, 0, 1, 1),
		(drawing, 6435, 6435, 0, 0, 0, 0, 1, 1),
		(drawing, 6434, 6434, 0, 0, 0, 0, 1, 1),
		(drawing, 6433, 6433, 0, 0, 0, 0, 1, 1),
		(drawing, 6432, 6432, 0, 0, 0, 0, 1, 1),
		(drawing, 6431, 6431, 0, 0, 0, 0, 1, 1),
		(drawing, 6430, 6430, 0, 0, 0, 0, 1, 1),
		(drawing, 6429, 6429, 0, 0, 0, 0, 1, 1),
		(drawing, 6428, 6428, 0, 0, 0, 0, 1, 1),
		(drawing, 6427, 6427, 0, 0, 0, 0, 1, 1),
		(drawing, 6426, 6426, 0, 0, 0, 0, 1, 1),
		(drawing, 6425, 6425, 0, 0, 0, 0, 1, 1),
		(drawing, 6424, 6424, 0, 0, 0, 0, 1, 1),
		(drawing, 6423, 6423, 0, 0, 0, 0, 1, 1),
		(drawing, 6422, 6422, 0, 0, 0, 0, 1, 1),
		(drawing, 6421, 6421, 0, 0, 0, 0, 1, 1),
		(drawing, 6420, 6420, 0, 0, 0, 0, 1, 1),
		(drawing, 6419, 6419, 0, 0, 0, 0, 1, 1),
		(drawing, 6418, 6418, 0, 0, 0, 0, 1, 1),
		(drawing, 6417, 6417, 0, 0, 0, 0, 1, 1),
		(drawing, 6416, 6416, 0, 0, 0, 0, 1, 1),
		(drawing, 6415, 6415, 0, 0, 0, 0, 1, 1),
		(drawing, 6414, 6414, 0, 0, 0, 0, 1, 1),
		(drawing, 6413, 6413, 0, 0, 0, 0, 1, 1),
		(drawing, 6412, 6412, 0, 0, 0, 0, 1, 1),
		(drawing, 6411, 6411, 0, 0, 0, 0, 1, 1),
		(drawing, 6410, 6410, 0, 0, 0, 0, 1, 1),
		(drawing, 6409, 6409, 0, 0, 0, 0, 1, 1),
		(drawing, 6408, 6408, 0, 0, 0, 0, 1, 1),
		(drawing, 6407, 6407, 0, 0, 0, 0, 1, 1),
		(drawing, 6406, 6406, 0, 0, 0, 0, 1, 1),
		(drawing, 6405, 6405, 0, 0, 0, 0, 1, 1),
		(drawing, 6404, 6404, 0, 0, 0, 0, 1, 1),
		(drawing, 6403, 6403, 0, 0, 0, 0, 1, 1),
		(drawing, 6402, 6402, 0, 0, 0, 0, 1, 1),
		(drawing, 6401, 6401, 0, 0, 0, 0, 1, 1),
		(drawing, 6400, 6400, 0, 0, 0, 0, 1, 1),
		(drawing, 6399, 6399, 0, 0, 0, 0, 1, 1),
		(drawing, 6398, 6398, 0, 0, 0, 0, 1, 1),
		(drawing, 6397, 6397, 0, 0, 0, 0, 1, 1),
		(drawing, 6396, 6396, 0, 0, 0, 0, 1, 1),
		(drawing, 6395, 6395, 0, 0, 0, 0, 1, 1),
		(drawing, 6394, 6394, 0, 0, 0, 0, 1, 1),
		(drawing, 6393, 6393, 0, 0, 0, 0, 1, 1),
		(drawing, 6392, 6392, 0, 0, 0, 0, 1, 1),
		(drawing, 6391, 6391, 0, 0, 0, 0, 1, 1),
		(drawing, 6390, 6390, 0, 0, 0, 0, 1, 1),
		(drawing, 6389, 6389, 0, 0, 0, 0, 1, 1),
		(drawing, 6388, 6388, 0, 0, 0, 0, 1, 1),
		(drawing, 6387, 6387, 0, 0, 0, 0, 1, 1),
		(drawing, 6386, 6386, 0, 0, 0, 0, 1, 1),
		(drawing, 6385, 6385, 0, 0, 0, 0, 1, 1),
		(drawing, 6384, 6384, 0, 0, 0, 0, 1, 1),
		(drawing, 6383, 6383, 0, 0, 0, 0, 1, 1),
		(drawing, 6382, 6382, 0, 0, 0, 0, 1, 1),
		(drawing, 6381, 6381, 0, 0, 0, 0, 1, 1),
		(drawing, 6380, 6380, 0, 0, 0, 0, 1, 1),
		(drawing, 6379, 6379, 0, 0, 0, 0, 1, 1),
		(drawing, 6378, 6378, 0, 0, 0, 0, 1, 1),
		(drawing, 6377, 6377, 0, 0, 0, 0, 1, 1),
		(drawing, 6376, 6376, 0, 0, 0, 0, 1, 1),
		(drawing, 6375, 6375, 0, 0, 0, 0, 1, 1),
		(drawing, 6374, 6374, 0, 0, 0, 0, 1, 1),
		(drawing, 6373, 6373, 0, 0, 0, 0, 1, 1),
		(drawing, 6372, 6372, 0, 0, 0, 0, 1, 1),
		(drawing, 6371, 6371, 0, 0, 0, 0, 1, 1),
		(drawing, 6370, 6370, 0, 0, 0, 0, 1, 1),
		(drawing, 6369, 6369, 0, 0, 0, 0, 1, 1),
		(drawing, 6368, 6368, 0, 0, 0, 0, 1, 1),
		(drawing, 6367, 6367, 0, 0, 0, 0, 1, 1),
		(drawing, 6366, 6366, 0, 0, 0, 0, 1, 1),
		(drawing, 6365, 6365, 0, 0, 0, 0, 1, 1),
		(drawing, 6364, 6364, 0, 0, 0, 0, 1, 1),
		(drawing, 6363, 6363, 0, 0, 0, 0, 1, 1),
		(drawing, 6362, 6362, 0, 0, 0, 0, 1, 1),
		(drawing, 6361, 6361, 0, 0, 0, 0, 1, 1),
		(drawing, 6360, 6360, 0, 0, 0, 0, 1, 1),
		(drawing, 6359, 6359, 0, 0, 0, 0, 1, 1),
		(drawing, 6358, 6358, 0, 0, 0, 0, 1, 1),
		(drawing, 6357, 6357, 0, 0, 0, 0, 1, 1),
		(drawing, 6356, 6356, 0, 0, 0, 0, 1, 1),
		(drawing, 6355, 6355, 0, 0, 0, 0, 1, 1),
		(drawing, 6354, 6354, 0, 0, 0, 0, 1, 1),
		(drawing, 6353, 6353, 0, 0, 0, 0, 1, 1),
		(drawing, 6352, 6352, 0, 0, 0, 0, 1, 1),
		(drawing, 6351, 6351, 0, 0, 0, 0, 1, 1),
		(drawing, 6350, 6350, 0, 0, 0, 0, 1, 1),
		(drawing, 6349, 6349, 0, 0, 0, 0, 1, 1),
		(drawing, 6348, 6348, 0, 0, 0, 0, 1, 1),
		(drawing, 6347, 6347, 0, 0, 0, 0, 1, 1),
		(drawing, 6346, 6346, 0, 0, 0, 0, 1, 1),
		(drawing, 6345, 6345, 0, 0, 0, 0, 1, 1),
		(drawing, 6344, 6344, 0, 0, 0, 0, 1, 1),
		(drawing, 6343, 6343, 0, 0, 0, 0, 1, 1),
		(drawing, 6342, 6342, 0, 0, 0, 0, 1, 1),
		(drawing, 6341, 6341, 0, 0, 0, 0, 1, 1),
		(drawing, 6340, 6340, 0, 0, 0, 0, 1, 1),
		(drawing, 6339, 6339, 0, 0, 0, 0, 1, 1),
		(drawing, 6338, 6338, 0, 0, 0, 0, 1, 1),
		(drawing, 6337, 6337, 0, 0, 0, 0, 1, 1),
		(drawing, 6336, 6336, 0, 0, 0, 0, 1, 1),
		(drawing, 6335, 6335, 0, 0, 0, 0, 1, 1),
		(drawing, 6334, 6334, 0, 0, 0, 0, 1, 1),
		(drawing, 6333, 6333, 0, 0, 0, 0, 1, 1),
		(drawing, 6332, 6332, 0, 0, 0, 0, 1, 1),
		(drawing, 6331, 6331, 0, 0, 0, 0, 1, 1),
		(drawing, 6330, 6330, 0, 0, 0, 0, 1, 1),
		(drawing, 6329, 6329, 0, 0, 0, 0, 1, 1),
		(drawing, 6328, 6328, 0, 0, 0, 0, 1, 1),
		(drawing, 6327, 6327, 0, 0, 0, 0, 1, 1),
		(drawing, 6326, 6326, 0, 0, 0, 0, 1, 1),
		(drawing, 6325, 6325, 0, 0, 0, 0, 1, 1),
		(drawing, 6324, 6324, 0, 0, 0, 0, 1, 1),
		(drawing, 6323, 6323, 0, 0, 0, 0, 1, 1),
		(drawing, 6322, 6322, 0, 0, 0, 0, 1, 1),
		(drawing, 6321, 6321, 0, 0, 0, 0, 1, 1),
		(drawing, 6320, 6320, 0, 0, 0, 0, 1, 1),
		(drawing, 6319, 6319, 0, 0, 0, 0, 1, 1),
		(drawing, 6318, 6318, 0, 0, 0, 0, 1, 1),
		(drawing, 6317, 6317, 0, 0, 0, 0, 1, 1),
		(drawing, 6316, 6316, 0, 0, 0, 0, 1, 1),
		(drawing, 6315, 6315, 0, 0, 0, 0, 1, 1),
		(drawing, 6314, 6314, 0, 0, 0, 0, 1, 1),
		(drawing, 6313, 6313, 0, 0, 0, 0, 1, 1),
		(drawing, 6312, 6312, 0, 0, 0, 0, 1, 1),
		(drawing, 6311, 6311, 0, 0, 0, 0, 1, 1),
		(drawing, 6310, 6310, 0, 0, 0, 0, 1, 1),
		(drawing, 6309, 6309, 0, 0, 0, 0, 1, 1),
		(drawing, 6308, 6308, 0, 0, 0, 0, 1, 1),
		(drawing, 6307, 6307, 0, 0, 0, 0, 1, 1),
		(drawing, 6306, 6306, 0, 0, 0, 0, 1, 1),
		(drawing, 6305, 6305, 0, 0, 0, 0, 1, 1),
		(drawing, 6304, 6304, 0, 0, 0, 0, 1, 1),
		(drawing, 6303, 6303, 0, 0, 0, 0, 1, 1),
		(drawing, 6302, 6302, 0, 0, 0, 0, 1, 1),
		(drawing, 6301, 6301, 0, 0, 0, 0, 1, 1),
		(drawing, 6300, 6300, 0, 0, 0, 0, 1, 1),
		(drawing, 6299, 6299, 0, 0, 0, 0, 1, 1),
		(drawing, 6298, 6298, 0, 0, 0, 0, 1, 1),
		(drawing, 6297, 6297, 0, 0, 0, 0, 1, 1),
		(drawing, 6296, 6296, 0, 0, 0, 0, 1, 1),
		(drawing, 6295, 6295, 0, 0, 0, 0, 1, 1),
		(drawing, 6294, 6294, 0, 0, 0, 0, 1, 1),
		(drawing, 6293, 6293, 0, 0, 0, 0, 1, 1),
		(drawing, 6292, 6292, 0, 0, 0, 0, 1, 1),
		(drawing, 6291, 6291, 0, 0, 0, 0, 1, 1),
		(drawing, 6290, 6290, 0, 0, 0, 0, 1, 1),
		(drawing, 6289, 6289, 0, 0, 0, 0, 1, 1),
		(drawing, 6288, 6288, 0, 0, 0, 0, 1, 1),
		(drawing, 6287, 6287, 0, 0, 0, 0, 1, 1),
		(drawing, 6286, 6286, 0, 0, 0, 0, 1, 1),
		(drawing, 6285, 6285, 0, 0, 0, 0, 1, 1),
		(drawing, 6284, 6284, 0, 0, 0, 0, 1, 1),
		(drawing, 6283, 6283, 0, 0, 0, 0, 1, 1),
		(drawing, 6282, 6282, 0, 0, 0, 0, 1, 1),
		(drawing, 6281, 6281, 0, 0, 0, 0, 1, 1),
		(drawing, 6280, 6280, 0, 0, 0, 0, 1, 1),
		(drawing, 6279, 6279, 0, 0, 0, 0, 1, 1),
		(drawing, 6278, 6278, 0, 0, 0, 0, 1, 1),
		(drawing, 6277, 6277, 0, 0, 0, 0, 1, 1),
		(drawing, 6276, 6276, 0, 0, 0, 0, 1, 1),
		(drawing, 6275, 6275, 0, 0, 0, 0, 1, 1),
		(drawing, 6274, 6274, 0, 0, 0, 0, 1, 1),
		(drawing, 6273, 6273, 0, 0, 0, 0, 1, 1),
		(drawing, 6272, 6272, 0, 0, 0, 0, 1, 1),
		(drawing, 6271, 6271, 0, 0, 0, 0, 1, 1),
		(drawing, 6270, 6270, 0, 0, 0, 0, 1, 1),
		(drawing, 6269, 6269, 0, 0, 0, 0, 1, 1),
		(drawing, 6268, 6268, 0, 0, 0, 0, 1, 1),
		(drawing, 6267, 6267, 0, 0, 0, 0, 1, 1),
		(drawing, 6266, 6266, 0, 0, 0, 0, 1, 1),
		(drawing, 6265, 6265, 0, 0, 0, 0, 1, 1),
		(drawing, 6264, 6264, 0, 0, 0, 0, 1, 1),
		(drawing, 6263, 6263, 0, 0, 0, 0, 1, 1),
		(drawing, 6262, 6262, 0, 0, 0, 0, 1, 1),
		(drawing, 6261, 6261, 0, 0, 0, 0, 1, 1),
		(drawing, 6260, 6260, 0, 0, 0, 0, 1, 1),
		(drawing, 6259, 6259, 0, 0, 0, 0, 1, 1),
		(drawing, 6258, 6258, 0, 0, 0, 0, 1, 1),
		(drawing, 6257, 6257, 0, 0, 0, 0, 1, 1),
		(drawing, 6256, 6256, 0, 0, 0, 0, 1, 1),
		(drawing, 6255, 6255, 0, 0, 0, 0, 1, 1),
		(drawing, 6254, 6254, 0, 0, 0, 0, 1, 1),
		(drawing, 6253, 6253, 0, 0, 0, 0, 1, 1),
		(drawing, 6252, 6252, 0, 0, 0, 0, 1, 1),
		(drawing, 6251, 6251, 0, 0, 0, 0, 1, 1),
		(drawing, 6250, 6250, 0, 0, 0, 0, 1, 1),
		(drawing, 6249, 6249, 0, 0, 0, 0, 1, 1),
		(drawing, 6248, 6248, 0, 0, 0, 0, 1, 1),
		(drawing, 6247, 6247, 0, 0, 0, 0, 1, 1),
		(drawing, 6246, 6246, 0, 0, 0, 0, 1, 1),
		(drawing, 6245, 6245, 0, 0, 0, 0, 1, 1),
		(drawing, 6244, 6244, 0, 0, 0, 0, 1, 1),
		(drawing, 6243, 6243, 0, 0, 0, 0, 1, 1),
		(drawing, 6242, 6242, 0, 0, 0, 0, 1, 1),
		(drawing, 6241, 6241, 0, 0, 0, 0, 1, 1),
		(drawing, 6240, 6240, 0, 0, 0, 0, 1, 1),
		(drawing, 6239, 6239, 0, 0, 0, 0, 1, 1),
		(drawing, 6238, 6238, 0, 0, 0, 0, 1, 1),
		(drawing, 6237, 6237, 0, 0, 0, 0, 1, 1),
		(drawing, 6236, 6236, 0, 0, 0, 0, 1, 1),
		(drawing, 6235, 6235, 0, 0, 0, 0, 1, 1),
		(drawing, 6234, 6234, 0, 0, 0, 0, 1, 1),
		(drawing, 6233, 6233, 0, 0, 0, 0, 1, 1),
		(drawing, 6232, 6232, 0, 0, 0, 0, 1, 1),
		(drawing, 6231, 6231, 0, 0, 0, 0, 1, 1),
		(drawing, 6230, 6230, 0, 0, 0, 0, 1, 1),
		(drawing, 6229, 6229, 0, 0, 0, 0, 1, 1),
		(drawing, 6228, 6228, 0, 0, 0, 0, 1, 1),
		(drawing, 6227, 6227, 0, 0, 0, 0, 1, 1),
		(drawing, 6226, 6226, 0, 0, 0, 0, 1, 1),
		(drawing, 6225, 6225, 0, 0, 0, 0, 1, 1),
		(drawing, 6224, 6224, 0, 0, 0, 0, 1, 1),
		(drawing, 6223, 6223, 0, 0, 0, 0, 1, 1),
		(drawing, 6222, 6222, 0, 0, 0, 0, 1, 1),
		(drawing, 6221, 6221, 0, 0, 0, 0, 1, 1),
		(drawing, 6220, 6220, 0, 0, 0, 0, 1, 1),
		(drawing, 6219, 6219, 0, 0, 0, 0, 1, 1),
		(drawing, 6218, 6218, 0, 0, 0, 0, 1, 1),
		(drawing, 6217, 6217, 0, 0, 0, 0, 1, 1),
		(drawing, 6216, 6216, 0, 0, 0, 0, 1, 1),
		(drawing, 6215, 6215, 0, 0, 0, 0, 1, 1),
		(drawing, 6214, 6214, 0, 0, 0, 0, 1, 1),
		(drawing, 6213, 6213, 0, 0, 0, 0, 1, 1),
		(drawing, 6212, 6212, 0, 0, 0, 0, 1, 1),
		(drawing, 6211, 6211, 0, 0, 0, 0, 1, 1),
		(drawing, 6210, 6210, 0, 0, 0, 0, 1, 1),
		(drawing, 6209, 6209, 0, 0, 0, 0, 1, 1),
		(drawing, 6208, 6208, 0, 0, 0, 0, 1, 1),
		(drawing, 6207, 6207, 0, 0, 0, 0, 1, 1),
		(drawing, 6206, 6206, 0, 0, 0, 0, 1, 1),
		(drawing, 6205, 6205, 0, 0, 0, 0, 1, 1),
		(drawing, 6204, 6204, 0, 0, 0, 0, 1, 1),
		(drawing, 6203, 6203, 0, 0, 0, 0, 1, 1),
		(drawing, 6202, 6202, 0, 0, 0, 0, 1, 1),
		(drawing, 6201, 6201, 0, 0, 0, 0, 1, 1),
		(drawing, 6200, 6200, 0, 0, 0, 0, 1, 1),
		(drawing, 6199, 6199, 0, 0, 0, 0, 1, 1),
		(drawing, 6198, 6198, 0, 0, 0, 0, 1, 1),
		(drawing, 6197, 6197, 0, 0, 0, 0, 1, 1),
		(drawing, 6196, 6196, 0, 0, 0, 0, 1, 1),
		(drawing, 6195, 6195, 0, 0, 0, 0, 1, 1),
		(drawing, 6194, 6194, 0, 0, 0, 0, 1, 1),
		(drawing, 6193, 6193, 0, 0, 0, 0, 1, 1),
		(drawing, 6192, 6192, 0, 0, 0, 0, 1, 1),
		(drawing, 6191, 6191, 0, 0, 0, 0, 1, 1),
		(drawing, 6190, 6190, 0, 0, 0, 0, 1, 1),
		(drawing, 6189, 6189, 0, 0, 0, 0, 1, 1),
		(drawing, 6188, 6188, 0, 0, 0, 0, 1, 1),
		(drawing, 6187, 6187, 0, 0, 0, 0, 1, 1),
		(drawing, 6186, 6186, 0, 0, 0, 0, 1, 1),
		(drawing, 6185, 6185, 0, 0, 0, 0, 1, 1),
		(drawing, 6184, 6184, 0, 0, 0, 0, 1, 1),
		(drawing, 6183, 6183, 0, 0, 0, 0, 1, 1),
		(drawing, 6182, 6182, 0, 0, 0, 0, 1, 1),
		(drawing, 6181, 6181, 0, 0, 0, 0, 1, 1),
		(drawing, 6180, 6180, 0, 0, 0, 0, 1, 1),
		(drawing, 6179, 6179, 0, 0, 0, 0, 1, 1),
		(drawing, 6178, 6178, 0, 0, 0, 0, 1, 1),
		(drawing, 6177, 6177, 0, 0, 0, 0, 1, 1),
		(drawing, 6176, 6176, 0, 0, 0, 0, 1, 1),
		(drawing, 6175, 6175, 0, 0, 0, 0, 1, 1),
		(drawing, 6174, 6174, 0, 0, 0, 0, 1, 1),
		(drawing, 6173, 6173, 0, 0, 0, 0, 1, 1),
		(drawing, 6172, 6172, 0, 0, 0, 0, 1, 1),
		(drawing, 6171, 6171, 0, 0, 0, 0, 1, 1),
		(drawing, 6170, 6170, 0, 0, 0, 0, 1, 1),
		(drawing, 6169, 6169, 0, 0, 0, 0, 1, 1),
		(drawing, 6168, 6168, 0, 0, 0, 0, 1, 1),
		(drawing, 6167, 6167, 0, 0, 0, 0, 1, 1),
		(drawing, 6166, 6166, 0, 0, 0, 0, 1, 1),
		(drawing, 6165, 6165, 0, 0, 0, 0, 1, 1),
		(drawing, 6164, 6164, 0, 0, 0, 0, 1, 1),
		(drawing, 6163, 6163, 0, 0, 0, 0, 1, 1),
		(drawing, 6162, 6162, 0, 0, 0, 0, 1, 1),
		(drawing, 6161, 6161, 0, 0, 0, 0, 1, 1),
		(drawing, 6160, 6160, 0, 0, 0, 0, 1, 1),
		(drawing, 6159, 6159, 0, 0, 0, 0, 1, 1),
		(drawing, 6158, 6158, 0, 0, 0, 0, 1, 1),
		(drawing, 6157, 6157, 0, 0, 0, 0, 1, 1),
		(drawing, 6156, 6156, 0, 0, 0, 0, 1, 1),
		(drawing, 6155, 6155, 0, 0, 0, 0, 1, 1),
		(drawing, 6154, 6154, 0, 0, 0, 0, 1, 1),
		(drawing, 6153, 6153, 0, 0, 0, 0, 1, 1),
		(drawing, 6152, 6152, 0, 0, 0, 0, 1, 1),
		(drawing, 6151, 6151, 0, 0, 0, 0, 1, 1),
		(drawing, 6150, 6150, 0, 0, 0, 0, 1, 1),
		(drawing, 6149, 6149, 0, 0, 0, 0, 1, 1),
		(drawing, 6148, 6148, 0, 0, 0, 0, 1, 1),
		(drawing, 6147, 6147, 0, 0, 0, 0, 1, 1),
		(drawing, 6146, 6146, 0, 0, 0, 0, 1, 1),
		(drawing, 6145, 6145, 0, 0, 0, 0, 1, 1),
		(drawing, 6144, 6144, 0, 0, 0, 0, 1, 1),
		(drawing, 6143, 6143, 0, 0, 0, 0, 1, 1),
		(drawing, 6142, 6142, 0, 0, 0, 0, 1, 1),
		(drawing, 6141, 6141, 0, 0, 0, 0, 1, 1),
		(drawing, 6140, 6140, 0, 0, 0, 0, 1, 1),
		(drawing, 6139, 6139, 0, 0, 0, 0, 1, 1),
		(drawing, 6138, 6138, 0, 0, 0, 0, 1, 1),
		(drawing, 6137, 6137, 0, 0, 0, 0, 1, 1),
		(drawing, 6136, 6136, 0, 0, 0, 0, 1, 1),
		(drawing, 6135, 6135, 0, 0, 0, 0, 1, 1),
		(drawing, 6134, 6134, 0, 0, 0, 0, 1, 1),
		(drawing, 6133, 6133, 0, 0, 0, 0, 1, 1),
		(drawing, 6132, 6132, 0, 0, 0, 0, 1, 1),
		(drawing, 6131, 6131, 0, 0, 0, 0, 1, 1),
		(drawing, 6130, 6130, 0, 0, 0, 0, 1, 1),
		(drawing, 6129, 6129, 0, 0, 0, 0, 1, 1),
		(drawing, 6128, 6128, 0, 0, 0, 0, 1, 1),
		(drawing, 6127, 6127, 0, 0, 0, 0, 1, 1),
		(drawing, 6126, 6126, 0, 0, 0, 0, 1, 1),
		(drawing, 6125, 6125, 0, 0, 0, 0, 1, 1),
		(drawing, 6124, 6124, 0, 0, 0, 0, 1, 1),
		(drawing, 6123, 6123, 0, 0, 0, 0, 1, 1),
		(drawing, 6122, 6122, 0, 0, 0, 0, 1, 1),
		(drawing, 6121, 6121, 0, 0, 0, 0, 1, 1),
		(drawing, 6120, 6120, 0, 0, 0, 0, 1, 1),
		(drawing, 6119, 6119, 0, 0, 0, 0, 1, 1),
		(drawing, 6118, 6118, 0, 0, 0, 0, 1, 1),
		(drawing, 6117, 6117, 0, 0, 0, 0, 1, 1),
		(drawing, 6116, 6116, 0, 0, 0, 0, 1, 1),
		(drawing, 6115, 6115, 0, 0, 0, 0, 1, 1),
		(drawing, 6114, 6114, 0, 0, 0, 0, 1, 1),
		(drawing, 6113, 6113, 0, 0, 0, 0, 1, 1),
		(drawing, 6112, 6112, 0, 0, 0, 0, 1, 1),
		(drawing, 6111, 6111, 0, 0, 0, 0, 1, 1),
		(drawing, 6110, 6110, 0, 0, 0, 0, 1, 1),
		(drawing, 6109, 6109, 0, 0, 0, 0, 1, 1),
		(drawing, 6108, 6108, 0, 0, 0, 0, 1, 1),
		(drawing, 6107, 6107, 0, 0, 0, 0, 1, 1),
		(drawing, 6106, 6106, 0, 0, 0, 0, 1, 1),
		(drawing, 6105, 6105, 0, 0, 0, 0, 1, 1),
		(drawing, 6104, 6104, 0, 0, 0, 0, 1, 1),
		(drawing, 6103, 6103, 0, 0, 0, 0, 1, 1),
		(drawing, 6102, 6102, 0, 0, 0, 0, 1, 1),
		(drawing, 6101, 6101, 0, 0, 0, 0, 1, 1),
		(drawing, 6100, 6100, 0, 0, 0, 0, 1, 1),
		(drawing, 6099, 6099, 0, 0, 0, 0, 1, 1),
		(drawing, 6098, 6098, 0, 0, 0, 0, 1, 1),
		(drawing, 6097, 6097, 0, 0, 0, 0, 1, 1),
		(drawing, 6096, 6096, 0, 0, 0, 0, 1, 1),
		(drawing, 6095, 6095, 0, 0, 0, 0, 1, 1),
		(drawing, 6094, 6094, 0, 0, 0, 0, 1, 1),
		(drawing, 6093, 6093, 0, 0, 0, 0, 1, 1),
		(drawing, 6092, 6092, 0, 0, 0, 0, 1, 1),
		(drawing, 6091, 6091, 0, 0, 0, 0, 1, 1),
		(drawing, 6090, 6090, 0, 0, 0, 0, 1, 1),
		(drawing, 6089, 6089, 0, 0, 0, 0, 1, 1),
		(drawing, 6088, 6088, 0, 0, 0, 0, 1, 1),
		(drawing, 6087, 6087, 0, 0, 0, 0, 1, 1),
		(drawing, 6086, 6086, 0, 0, 0, 0, 1, 1),
		(drawing, 6085, 6085, 0, 0, 0, 0, 1, 1),
		(drawing, 6084, 6084, 0, 0, 0, 0, 1, 1),
		(drawing, 6083, 6083, 0, 0, 0, 0, 1, 1),
		(drawing, 6082, 6082, 0, 0, 0, 0, 1, 1),
		(drawing, 6081, 6081, 0, 0, 0, 0, 1, 1),
		(drawing, 6080, 6080, 0, 0, 0, 0, 1, 1),
		(drawing, 6079, 6079, 0, 0, 0, 0, 1, 1),
		(drawing, 6078, 6078, 0, 0, 0, 0, 1, 1),
		(drawing, 6077, 6077, 0, 0, 0, 0, 1, 1),
		(drawing, 6076, 6076, 0, 0, 0, 0, 1, 1),
		(drawing, 6075, 6075, 0, 0, 0, 0, 1, 1),
		(drawing, 6074, 6074, 0, 0, 0, 0, 1, 1),
		(drawing, 6073, 6073, 0, 0, 0, 0, 1, 1),
		(drawing, 6072, 6072, 0, 0, 0, 0, 1, 1),
		(drawing, 6071, 6071, 0, 0, 0, 0, 1, 1),
		(drawing, 6070, 6070, 0, 0, 0, 0, 1, 1),
		(drawing, 6069, 6069, 0, 0, 0, 0, 1, 1),
		(drawing, 6068, 6068, 0, 0, 0, 0, 1, 1),
		(drawing, 6067, 6067, 0, 0, 0, 0, 1, 1),
		(drawing, 6066, 6066, 0, 0, 0, 0, 1, 1),
		(drawing, 6065, 6065, 0, 0, 0, 0, 1, 1),
		(drawing, 6064, 6064, 0, 0, 0, 0, 1, 1),
		(drawing, 6063, 6063, 0, 0, 0, 0, 1, 1),
		(drawing, 6062, 6062, 0, 0, 0, 0, 1, 1),
		(drawing, 6061, 6061, 0, 0, 0, 0, 1, 1),
		(drawing, 6060, 6060, 0, 0, 0, 0, 1, 1),
		(drawing, 6059, 6059, 0, 0, 0, 0, 1, 1),
		(drawing, 6058, 6058, 0, 0, 0, 0, 1, 1),
		(drawing, 6057, 6057, 0, 0, 0, 0, 1, 1),
		(drawing, 6056, 6056, 0, 0, 0, 0, 1, 1),
		(drawing, 6055, 6055, 0, 0, 0, 0, 1, 1),
		(drawing, 6054, 6054, 0, 0, 0, 0, 1, 1),
		(drawing, 6053, 6053, 0, 0, 0, 0, 1, 1),
		(drawing, 6052, 6052, 0, 0, 0, 0, 1, 1),
		(drawing, 6051, 6051, 0, 0, 0, 0, 1, 1),
		(drawing, 6050, 6050, 0, 0, 0, 0, 1, 1),
		(drawing, 6049, 6049, 0, 0, 0, 0, 1, 1),
		(drawing, 6048, 6048, 0, 0, 0, 0, 1, 1),
		(drawing, 6047, 6047, 0, 0, 0, 0, 1, 1),
		(drawing, 6046, 6046, 0, 0, 0, 0, 1, 1),
		(drawing, 6045, 6045, 0, 0, 0, 0, 1, 1),
		(drawing, 6044, 6044, 0, 0, 0, 0, 1, 1),
		(drawing, 6043, 6043, 0, 0, 0, 0, 1, 1),
		(drawing, 6042, 6042, 0, 0, 0, 0, 1, 1),
		(drawing, 6041, 6041, 0, 0, 0, 0, 1, 1),
		(drawing, 6040, 6040, 0, 0, 0, 0, 1, 1),
		(drawing, 6039, 6039, 0, 0, 0, 0, 1, 1),
		(drawing, 6038, 6038, 0, 0, 0, 0, 1, 1),
		(drawing, 6037, 6037, 0, 0, 0, 0, 1, 1),
		(drawing, 6036, 6036, 0, 0, 0, 0, 1, 1),
		(drawing, 6035, 6035, 0, 0, 0, 0, 1, 1),
		(drawing, 6034, 6034, 0, 0, 0, 0, 1, 1),
		(drawing, 6033, 6033, 0, 0, 0, 0, 1, 1),
		(drawing, 6032, 6032, 0, 0, 0, 0, 1, 1),
		(drawing, 6031, 6031, 0, 0, 0, 0, 1, 1),
		(drawing, 6030, 6030, 0, 0, 0, 0, 1, 1),
		(drawing, 6029, 6029, 0, 0, 0, 0, 1, 1),
		(drawing, 6028, 6028, 0, 0, 0, 0, 1, 1),
		(drawing, 6027, 6027, 0, 0, 0, 0, 1, 1),
		(drawing, 6026, 6026, 0, 0, 0, 0, 1, 1),
		(drawing, 6025, 6025, 0, 0, 0, 0, 1, 1),
		(drawing, 6024, 6024, 0, 0, 0, 0, 1, 1),
		(drawing, 6023, 6023, 0, 0, 0, 0, 1, 1),
		(drawing, 6022, 6022, 0, 0, 0, 0, 1, 1),
		(drawing, 6021, 6021, 0, 0, 0, 0, 1, 1),
		(drawing, 6020, 6020, 0, 0, 0, 0, 1, 1),
		(drawing, 6019, 6019, 0, 0, 0, 0, 1, 1),
		(drawing, 6018, 6018, 0, 0, 0, 0, 1, 1),
		(drawing, 6017, 6017, 0, 0, 0, 0, 1, 1),
		(drawing, 6016, 6016, 0, 0, 0, 0, 1, 1),
		(drawing, 6015, 6015, 0, 0, 0, 0, 1, 1),
		(drawing, 6014, 6014, 0, 0, 0, 0, 1, 1),
		(drawing, 6013, 6013, 0, 0, 0, 0, 1, 1),
		(drawing, 6012, 6012, 0, 0, 0, 0, 1, 1),
		(drawing, 6011, 6011, 0, 0, 0, 0, 1, 1),
		(drawing, 6010, 6010, 0, 0, 0, 0, 1, 1),
		(drawing, 6009, 6009, 0, 0, 0, 0, 1, 1),
		(drawing, 6008, 6008, 0, 0, 0, 0, 1, 1),
		(drawing, 6007, 6007, 0, 0, 0, 0, 1, 1),
		(drawing, 6006, 6006, 0, 0, 0, 0, 1, 1),
		(drawing, 6005, 6005, 0, 0, 0, 0, 1, 1),
		(drawing, 6004, 6004, 0, 0, 0, 0, 1, 1),
		(drawing, 6003, 6003, 0, 0, 0, 0, 1, 1),
		(drawing, 6002, 6002, 0, 0, 0, 0, 1, 1),
		(drawing, 6001, 6001, 0, 0, 0, 0, 1, 1),
		(drawing, 6000, 6000, 0, 0, 0, 0, 1, 1),
		(drawing, 5999, 5999, 0, 0, 0, 0, 1, 1),
		(drawing, 5998, 5998, 0, 0, 0, 0, 1, 1),
		(drawing, 5997, 5997, 0, 0, 0, 0, 1, 1),
		(drawing, 5996, 5996, 0, 0, 0, 0, 1, 1),
		(drawing, 5995, 5995, 0, 0, 0, 0, 1, 1),
		(drawing, 5994, 5994, 0, 0, 0, 0, 1, 1),
		(drawing, 5993, 5993, 0, 0, 0, 0, 1, 1),
		(drawing, 5992, 5992, 0, 0, 0, 0, 1, 1),
		(drawing, 5991, 5991, 0, 0, 0, 0, 1, 1),
		(drawing, 5990, 5990, 0, 0, 0, 0, 1, 1),
		(drawing, 5989, 5989, 0, 0, 0, 0, 1, 1),
		(drawing, 5988, 5988, 0, 0, 0, 0, 1, 1),
		(drawing, 5987, 5987, 0, 0, 0, 0, 1, 1),
		(drawing, 5986, 5986, 0, 0, 0, 0, 1, 1),
		(drawing, 5985, 5985, 0, 0, 0, 0, 1, 1),
		(drawing, 5984, 5984, 0, 0, 0, 0, 1, 1),
		(drawing, 5983, 5983, 0, 0, 0, 0, 1, 1),
		(drawing, 5982, 5982, 0, 0, 0, 0, 1, 1),
		(drawing, 5981, 5981, 0, 0, 0, 0, 1, 1),
		(drawing, 5980, 5980, 0, 0, 0, 0, 1, 1),
		(drawing, 5979, 5979, 0, 0, 0, 0, 1, 1),
		(drawing, 5978, 5978, 0, 0, 0, 0, 1, 1),
		(drawing, 5977, 5977, 0, 0, 0, 0, 1, 1),
		(drawing, 5976, 5976, 0, 0, 0, 0, 1, 1),
		(drawing, 5975, 5975, 0, 0, 0, 0, 1, 1),
		(drawing, 5974, 5974, 0, 0, 0, 0, 1, 1),
		(drawing, 5973, 5973, 0, 0, 0, 0, 1, 1),
		(drawing, 5972, 5972, 0, 0, 0, 0, 1, 1),
		(drawing, 5971, 5971, 0, 0, 0, 0, 1, 1),
		(drawing, 5970, 5970, 0, 0, 0, 0, 1, 1),
		(drawing, 5969, 5969, 0, 0, 0, 0, 1, 1),
		(drawing, 5968, 5968, 0, 0, 0, 0, 1, 1),
		(drawing, 5967, 5967, 0, 0, 0, 0, 1, 1),
		(drawing, 5966, 5966, 0, 0, 0, 0, 1, 1),
		(drawing, 5965, 5965, 0, 0, 0, 0, 1, 1),
		(drawing, 5964, 5964, 0, 0, 0, 0, 1, 1),
		(drawing, 5963, 5963, 0, 0, 0, 0, 1, 1),
		(drawing, 5962, 5962, 0, 0, 0, 0, 1, 1),
		(drawing, 5961, 5961, 0, 0, 0, 0, 1, 1),
		(drawing, 5960, 5960, 0, 0, 0, 0, 1, 1),
		(drawing, 5959, 5959, 0, 0, 0, 0, 1, 1),
		(drawing, 5958, 5958, 0, 0, 0, 0, 1, 1),
		(drawing, 5957, 5957, 0, 0, 0, 0, 1, 1),
		(drawing, 5956, 5956, 0, 0, 0, 0, 1, 1),
		(drawing, 5955, 5955, 0, 0, 0, 0, 1, 1),
		(drawing, 5954, 5954, 0, 0, 0, 0, 1, 1),
		(drawing, 5953, 5953, 0, 0, 0, 0, 1, 1),
		(drawing, 5952, 5952, 0, 0, 0, 0, 1, 1),
		(drawing, 5951, 5951, 0, 0, 0, 0, 1, 1),
		(drawing, 5950, 5950, 0, 0, 0, 0, 1, 1),
		(drawing, 5949, 5949, 0, 0, 0, 0, 1, 1),
		(drawing, 5948, 5948, 0, 0, 0, 0, 1, 1),
		(drawing, 5947, 5947, 0, 0, 0, 0, 1, 1),
		(drawing, 5946, 5946, 0, 0, 0, 0, 1, 1),
		(drawing, 5945, 5945, 0, 0, 0, 0, 1, 1),
		(drawing, 5944, 5944, 0, 0, 0, 0, 1, 1),
		(drawing, 5943, 5943, 0, 0, 0, 0, 1, 1),
		(drawing, 5942, 5942, 0, 0, 0, 0, 1, 1),
		(drawing, 5941, 5941, 0, 0, 0, 0, 1, 1),
		(drawing, 5940, 5940, 0, 0, 0, 0, 1, 1),
		(drawing, 5939, 5939, 0, 0, 0, 0, 1, 1),
		(drawing, 5938, 5938, 0, 0, 0, 0, 1, 1),
		(drawing, 5937, 5937, 0, 0, 0, 0, 1, 1),
		(drawing, 5936, 5936, 0, 0, 0, 0, 1, 1),
		(drawing, 5935, 5935, 0, 0, 0, 0, 1, 1),
		(drawing, 5934, 5934, 0, 0, 0, 0, 1, 1),
		(drawing, 5933, 5933, 0, 0, 0, 0, 1, 1),
		(drawing, 5932, 5932, 0, 0, 0, 0, 1, 1),
		(drawing, 5931, 5931, 0, 0, 0, 0, 1, 1),
		(drawing, 5930, 5930, 0, 0, 0, 0, 1, 1),
		(drawing, 5929, 5929, 0, 0, 0, 0, 1, 1),
		(drawing, 5928, 5928, 0, 0, 0, 0, 1, 1),
		(drawing, 5927, 5927, 0, 0, 0, 0, 1, 1),
		(drawing, 5926, 5926, 0, 0, 0, 0, 1, 1),
		(drawing, 5925, 5925, 0, 0, 0, 0, 1, 1),
		(drawing, 5924, 5924, 0, 0, 0, 0, 1, 1),
		(drawing, 5923, 5923, 0, 0, 0, 0, 1, 1),
		(drawing, 5922, 5922, 0, 0, 0, 0, 1, 1),
		(drawing, 5921, 5921, 0, 0, 0, 0, 1, 1),
		(drawing, 5920, 5920, 0, 0, 0, 0, 1, 1),
		(drawing, 5919, 5919, 0, 0, 0, 0, 1, 1),
		(drawing, 5918, 5918, 0, 0, 0, 0, 1, 1),
		(drawing, 5917, 5917, 0, 0, 0, 0, 1, 1),
		(drawing, 5916, 5916, 0, 0, 0, 0, 1, 1),
		(drawing, 5915, 5915, 0, 0, 0, 0, 1, 1),
		(drawing, 5914, 5914, 0, 0, 0, 0, 1, 1),
		(drawing, 5913, 5913, 0, 0, 0, 0, 1, 1),
		(drawing, 5912, 5912, 0, 0, 0, 0, 1, 1),
		(drawing, 5911, 5911, 0, 0, 0, 0, 1, 1),
		(drawing, 5910, 5910, 0, 0, 0, 0, 1, 1),
		(drawing, 5909, 5909, 0, 0, 0, 0, 1, 1),
		(drawing, 5908, 5908, 0, 0, 0, 0, 1, 1),
		(drawing, 5907, 5907, 0, 0, 0, 0, 1, 1),
		(drawing, 5906, 5906, 0, 0, 0, 0, 1, 1),
		(drawing, 5905, 5905, 0, 0, 0, 0, 1, 1),
		(drawing, 5904, 5904, 0, 0, 0, 0, 1, 1),
		(drawing, 5903, 5903, 0, 0, 0, 0, 1, 1),
		(drawing, 5902, 5902, 0, 0, 0, 0, 1, 1),
		(drawing, 5901, 5901, 0, 0, 0, 0, 1, 1),
		(drawing, 5900, 5900, 0, 0, 0, 0, 1, 1),
		(drawing, 5899, 5899, 0, 0, 0, 0, 1, 1),
		(drawing, 5898, 5898, 0, 0, 0, 0, 1, 1),
		(drawing, 5897, 5897, 0, 0, 0, 0, 1, 1),
		(drawing, 5896, 5896, 0, 0, 0, 0, 1, 1),
		(drawing, 5895, 5895, 0, 0, 0, 0, 1, 1),
		(drawing, 5894, 5894, 0, 0, 0, 0, 1, 1),
		(drawing, 5893, 5893, 0, 0, 0, 0, 1, 1),
		(drawing, 5892, 5892, 0, 0, 0, 0, 1, 1),
		(drawing, 5891, 5891, 0, 0, 0, 0, 1, 1),
		(drawing, 5890, 5890, 0, 0, 0, 0, 1, 1),
		(drawing, 5889, 5889, 0, 0, 0, 0, 1, 1),
		(drawing, 5888, 5888, 0, 0, 0, 0, 1, 1),
		(drawing, 5887, 5887, 0, 0, 0, 0, 1, 1),
		(drawing, 5886, 5886, 0, 0, 0, 0, 1, 1),
		(drawing, 5885, 5885, 0, 0, 0, 0, 1, 1),
		(drawing, 5884, 5884, 0, 0, 0, 0, 1, 1),
		(drawing, 5883, 5883, 0, 0, 0, 0, 1, 1),
		(drawing, 5882, 5882, 0, 0, 0, 0, 1, 1),
		(drawing, 5881, 5881, 0, 0, 0, 0, 1, 1),
		(drawing, 5880, 5880, 0, 0, 0, 0, 1, 1),
		(drawing, 5879, 5879, 0, 0, 0, 0, 1, 1),
		(drawing, 5878, 5878, 0, 0, 0, 0, 1, 1),
		(drawing, 5877, 5877, 0, 0, 0, 0, 1, 1),
		(drawing, 5876, 5876, 0, 0, 0, 0, 1, 1),
		(drawing, 5875, 5875, 0, 0, 0, 0, 1, 1),
		(drawing, 5874, 5874, 0, 0, 0, 0, 1, 1),
		(drawing, 5873, 5873, 0, 0, 0, 0, 1, 1),
		(drawing, 5872, 5872, 0, 0, 0, 0, 1, 1),
		(drawing, 5871, 5871, 0, 0, 0, 0, 1, 1),
		(drawing, 5870, 5870, 0, 0, 0, 0, 1, 1),
		(drawing, 5869, 5869, 0, 0, 0, 0, 1, 1),
		(drawing, 5868, 5868, 0, 0, 0, 0, 1, 1),
		(drawing, 5867, 5867, 0, 0, 0, 0, 1, 1),
		(drawing, 5866, 5866, 0, 0, 0, 0, 1, 1),
		(drawing, 5865, 5865, 0, 0, 0, 0, 1, 1),
		(drawing, 5864, 5864, 0, 0, 0, 0, 1, 1),
		(drawing, 5863, 5863, 0, 0, 0, 0, 1, 1),
		(drawing, 5862, 5862, 0, 0, 0, 0, 1, 1),
		(drawing, 5861, 5861, 0, 0, 0, 0, 1, 1),
		(drawing, 5860, 5860, 0, 0, 0, 0, 1, 1),
		(drawing, 5859, 5859, 0, 0, 0, 0, 1, 1),
		(drawing, 5858, 5858, 0, 0, 0, 0, 1, 1),
		(drawing, 5857, 5857, 0, 0, 0, 0, 1, 1),
		(drawing, 5856, 5856, 0, 0, 0, 0, 1, 1),
		(drawing, 5855, 5855, 0, 0, 0, 0, 1, 1),
		(drawing, 5854, 5854, 0, 0, 0, 0, 1, 1),
		(drawing, 5853, 5853, 0, 0, 0, 0, 1, 1),
		(drawing, 5852, 5852, 0, 0, 0, 0, 1, 1),
		(drawing, 5851, 5851, 0, 0, 0, 0, 1, 1),
		(drawing, 5850, 5850, 0, 0, 0, 0, 1, 1),
		(drawing, 5849, 5849, 0, 0, 0, 0, 1, 1),
		(drawing, 5848, 5848, 0, 0, 0, 0, 1, 1),
		(drawing, 5847, 5847, 0, 0, 0, 0, 1, 1),
		(drawing, 5846, 5846, 0, 0, 0, 0, 1, 1),
		(drawing, 5845, 5845, 0, 0, 0, 0, 1, 1),
		(drawing, 5844, 5844, 0, 0, 0, 0, 1, 1),
		(drawing, 5843, 5843, 0, 0, 0, 0, 1, 1),
		(drawing, 5842, 5842, 0, 0, 0, 0, 1, 1),
		(drawing, 5841, 5841, 0, 0, 0, 0, 1, 1),
		(drawing, 5840, 5840, 0, 0, 0, 0, 1, 1),
		(drawing, 5839, 5839, 0, 0, 0, 0, 1, 1),
		(drawing, 5838, 5838, 0, 0, 0, 0, 1, 1),
		(drawing, 5837, 5837, 0, 0, 0, 0, 1, 1),
		(drawing, 5836, 5836, 0, 0, 0, 0, 1, 1),
		(drawing, 5835, 5835, 0, 0, 0, 0, 1, 1),
		(drawing, 5834, 5834, 0, 0, 0, 0, 1, 1),
		(drawing, 5833, 5833, 0, 0, 0, 0, 1, 1),
		(drawing, 5832, 5832, 0, 0, 0, 0, 1, 1),
		(drawing, 5831, 5831, 0, 0, 0, 0, 1, 1),
		(drawing, 5830, 5830, 0, 0, 0, 0, 1, 1),
		(drawing, 5829, 5829, 0, 0, 0, 0, 1, 1),
		(drawing, 5828, 5828, 0, 0, 0, 0, 1, 1),
		(drawing, 5827, 5827, 0, 0, 0, 0, 1, 1),
		(drawing, 5826, 5826, 0, 0, 0, 0, 1, 1),
		(drawing, 5825, 5825, 0, 0, 0, 0, 1, 1),
		(drawing, 5824, 5824, 0, 0, 0, 0, 1, 1),
		(drawing, 5823, 5823, 0, 0, 0, 0, 1, 1),
		(drawing, 5822, 5822, 0, 0, 0, 0, 1, 1),
		(drawing, 5821, 5821, 0, 0, 0, 0, 1, 1),
		(drawing, 5820, 5820, 0, 0, 0, 0, 1, 1),
		(drawing, 5819, 5819, 0, 0, 0, 0, 1, 1),
		(drawing, 5818, 5818, 0, 0, 0, 0, 1, 1),
		(drawing, 5817, 5817, 0, 0, 0, 0, 1, 1),
		(drawing, 5816, 5816, 0, 0, 0, 0, 1, 1),
		(drawing, 5815, 5815, 0, 0, 0, 0, 1, 1),
		(drawing, 5814, 5814, 0, 0, 0, 0, 1, 1),
		(drawing, 5813, 5813, 0, 0, 0, 0, 1, 1),
		(drawing, 5812, 5812, 0, 0, 0, 0, 1, 1),
		(drawing, 5811, 5811, 0, 0, 0, 0, 1, 1),
		(drawing, 5810, 5810, 0, 0, 0, 0, 1, 1),
		(drawing, 5809, 5809, 0, 0, 0, 0, 1, 1),
		(drawing, 5808, 5808, 0, 0, 0, 0, 1, 1),
		(drawing, 5807, 5807, 0, 0, 0, 0, 1, 1),
		(drawing, 5806, 5806, 0, 0, 0, 0, 1, 1),
		(drawing, 5805, 5805, 0, 0, 0, 0, 1, 1),
		(drawing, 5804, 5804, 0, 0, 0, 0, 1, 1),
		(drawing, 5803, 5803, 0, 0, 0, 0, 1, 1),
		(drawing, 5802, 5802, 0, 0, 0, 0, 1, 1),
		(drawing, 5801, 5801, 0, 0, 0, 0, 1, 1),
		(drawing, 5800, 5800, 0, 0, 0, 0, 1, 1),
		(drawing, 5799, 5799, 0, 0, 0, 0, 1, 1),
		(drawing, 5798, 5798, 0, 0, 0, 0, 1, 1),
		(drawing, 5797, 5797, 0, 0, 0, 0, 1, 1),
		(drawing, 5796, 5796, 0, 0, 0, 0, 1, 1),
		(drawing, 5795, 5795, 0, 0, 0, 0, 1, 1),
		(drawing, 5794, 5794, 0, 0, 0, 0, 1, 1),
		(drawing, 5793, 5793, 0, 0, 0, 0, 1, 1),
		(drawing, 5792, 5792, 0, 0, 0, 0, 1, 1),
		(drawing, 5791, 5791, 0, 0, 0, 0, 1, 1),
		(drawing, 5790, 5790, 0, 0, 0, 0, 1, 1),
		(drawing, 5789, 5789, 0, 0, 0, 0, 1, 1),
		(drawing, 5788, 5788, 0, 0, 0, 0, 1, 1),
		(drawing, 5787, 5787, 0, 0, 0, 0, 1, 1),
		(drawing, 5786, 5786, 0, 0, 0, 0, 1, 1),
		(drawing, 5785, 5785, 0, 0, 0, 0, 1, 1),
		(drawing, 5784, 5784, 0, 0, 0, 0, 1, 1),
		(drawing, 5783, 5783, 0, 0, 0, 0, 1, 1),
		(drawing, 5782, 5782, 0, 0, 0, 0, 1, 1),
		(drawing, 5781, 5781, 0, 0, 0, 0, 1, 1),
		(drawing, 5780, 5780, 0, 0, 0, 0, 1, 1),
		(drawing, 5779, 5779, 0, 0, 0, 0, 1, 1),
		(drawing, 5778, 5778, 0, 0, 0, 0, 1, 1),
		(drawing, 5777, 5777, 0, 0, 0, 0, 1, 1),
		(drawing, 5776, 5776, 0, 0, 0, 0, 1, 1),
		(drawing, 5775, 5775, 0, 0, 0, 0, 1, 1),
		(drawing, 5774, 5774, 0, 0, 0, 0, 1, 1),
		(drawing, 5773, 5773, 0, 0, 0, 0, 1, 1),
		(drawing, 5772, 5772, 0, 0, 0, 0, 1, 1),
		(drawing, 5771, 5771, 0, 0, 0, 0, 1, 1),
		(drawing, 5770, 5770, 0, 0, 0, 0, 1, 1),
		(drawing, 5769, 5769, 0, 0, 0, 0, 1, 1),
		(drawing, 5768, 5768, 0, 0, 0, 0, 1, 1),
		(drawing, 5767, 5767, 0, 0, 0, 0, 1, 1),
		(drawing, 5766, 5766, 0, 0, 0, 0, 1, 1),
		(drawing, 5765, 5765, 0, 0, 0, 0, 1, 1),
		(drawing, 5764, 5764, 0, 0, 0, 0, 1, 1),
		(drawing, 5763, 5763, 0, 0, 0, 0, 1, 1),
		(drawing, 5762, 5762, 0, 0, 0, 0, 1, 1),
		(drawing, 5761, 5761, 0, 0, 0, 0, 1, 1),
		(drawing, 5760, 5760, 0, 0, 0, 0, 1, 1),
		(drawing, 5759, 5759, 0, 0, 0, 0, 1, 1),
		(drawing, 5758, 5758, 0, 0, 0, 0, 1, 1),
		(drawing, 5757, 5757, 0, 0, 0, 0, 1, 1),
		(drawing, 5756, 5756, 0, 0, 0, 0, 1, 1),
		(drawing, 5755, 5755, 0, 0, 0, 0, 1, 1),
		(drawing, 5754, 5754, 0, 0, 0, 0, 1, 1),
		(drawing, 5753, 5753, 0, 0, 0, 0, 1, 1),
		(drawing, 5752, 5752, 0, 0, 0, 0, 1, 1),
		(drawing, 5751, 5751, 0, 0, 0, 0, 1, 1),
		(drawing, 5750, 5750, 0, 0, 0, 0, 1, 1),
		(drawing, 5749, 5749, 0, 0, 0, 0, 1, 1),
		(drawing, 5748, 5748, 0, 0, 0, 0, 1, 1),
		(drawing, 5747, 5747, 0, 0, 0, 0, 1, 1),
		(drawing, 5746, 5746, 0, 0, 0, 0, 1, 1),
		(drawing, 5745, 5745, 0, 0, 0, 0, 1, 1),
		(drawing, 5744, 5744, 0, 0, 0, 0, 1, 1),
		(drawing, 5743, 5743, 0, 0, 0, 0, 1, 1),
		(drawing, 5742, 5742, 0, 0, 0, 0, 1, 1),
		(drawing, 5741, 5741, 0, 0, 0, 0, 1, 1),
		(drawing, 5740, 5740, 0, 0, 0, 0, 1, 1),
		(drawing, 5739, 5739, 0, 0, 0, 0, 1, 1),
		(drawing, 5738, 5738, 0, 0, 0, 0, 1, 1),
		(drawing, 5737, 5737, 0, 0, 0, 0, 1, 1),
		(drawing, 5736, 5736, 0, 0, 0, 0, 1, 1),
		(drawing, 5735, 5735, 0, 0, 0, 0, 1, 1),
		(drawing, 5734, 5734, 0, 0, 0, 0, 1, 1),
		(drawing, 5733, 5733, 0, 0, 0, 0, 1, 1),
		(drawing, 5732, 5732, 0, 0, 0, 0, 1, 1),
		(drawing, 5731, 5731, 0, 0, 0, 0, 1, 1),
		(drawing, 5730, 5730, 0, 0, 0, 0, 1, 1),
		(drawing, 5729, 5729, 0, 0, 0, 0, 1, 1),
		(drawing, 5728, 5728, 0, 0, 0, 0, 1, 1),
		(drawing, 5727, 5727, 0, 0, 0, 0, 1, 1),
		(drawing, 5726, 5726, 0, 0, 0, 0, 1, 1),
		(drawing, 5725, 5725, 0, 0, 0, 0, 1, 1),
		(drawing, 5724, 5724, 0, 0, 0, 0, 1, 1),
		(drawing, 5723, 5723, 0, 0, 0, 0, 1, 1),
		(drawing, 5722, 5722, 0, 0, 0, 0, 1, 1),
		(drawing, 5721, 5721, 0, 0, 0, 0, 1, 1),
		(drawing, 5720, 5720, 0, 0, 0, 0, 1, 1),
		(drawing, 5719, 5719, 0, 0, 0, 0, 1, 1),
		(drawing, 5718, 5718, 0, 0, 0, 0, 1, 1),
		(drawing, 5717, 5717, 0, 0, 0, 0, 1, 1),
		(drawing, 5716, 5716, 0, 0, 0, 0, 1, 1),
		(drawing, 5715, 5715, 0, 0, 0, 0, 1, 1),
		(drawing, 5714, 5714, 0, 0, 0, 0, 1, 1),
		(drawing, 5713, 5713, 0, 0, 0, 0, 1, 1),
		(drawing, 5712, 5712, 0, 0, 0, 0, 1, 1),
		(drawing, 5711, 5711, 0, 0, 0, 0, 1, 1),
		(drawing, 5710, 5710, 0, 0, 0, 0, 1, 1),
		(drawing, 5709, 5709, 0, 0, 0, 0, 1, 1),
		(drawing, 5708, 5708, 0, 0, 0, 0, 1, 1),
		(drawing, 5707, 5707, 0, 0, 0, 0, 1, 1),
		(drawing, 5706, 5706, 0, 0, 0, 0, 1, 1),
		(drawing, 5705, 5705, 0, 0, 0, 0, 1, 1),
		(drawing, 5704, 5704, 0, 0, 0, 0, 1, 1),
		(drawing, 5703, 5703, 0, 0, 0, 0, 1, 1),
		(drawing, 5702, 5702, 0, 0, 0, 0, 1, 1),
		(drawing, 5701, 5701, 0, 0, 0, 0, 1, 1),
		(drawing, 5700, 5700, 0, 0, 0, 0, 1, 1),
		(drawing, 5699, 5699, 0, 0, 0, 0, 1, 1),
		(drawing, 5698, 5698, 0, 0, 0, 0, 1, 1),
		(drawing, 5697, 5697, 0, 0, 0, 0, 1, 1),
		(drawing, 5696, 5696, 0, 0, 0, 0, 1, 1),
		(drawing, 5695, 5695, 0, 0, 0, 0, 1, 1),
		(drawing, 5694, 5694, 0, 0, 0, 0, 1, 1),
		(drawing, 5693, 5693, 0, 0, 0, 0, 1, 1),
		(drawing, 5692, 5692, 0, 0, 0, 0, 1, 1),
		(drawing, 5691, 5691, 0, 0, 0, 0, 1, 1),
		(drawing, 5690, 5690, 0, 0, 0, 0, 1, 1),
		(drawing, 5689, 5689, 0, 0, 0, 0, 1, 1),
		(drawing, 5688, 5688, 0, 0, 0, 0, 1, 1),
		(drawing, 5687, 5687, 0, 0, 0, 0, 1, 1),
		(drawing, 5686, 5686, 0, 0, 0, 0, 1, 1),
		(drawing, 5685, 5685, 0, 0, 0, 0, 1, 1),
		(drawing, 5684, 5684, 0, 0, 0, 0, 1, 1),
		(drawing, 5683, 5683, 0, 0, 0, 0, 1, 1),
		(drawing, 5682, 5682, 0, 0, 0, 0, 1, 1),
		(drawing, 5681, 5681, 0, 0, 0, 0, 1, 1),
		(drawing, 5680, 5680, 0, 0, 0, 0, 1, 1),
		(drawing, 5679, 5679, 0, 0, 0, 0, 1, 1),
		(drawing, 5678, 5678, 0, 0, 0, 0, 1, 1),
		(drawing, 5677, 5677, 0, 0, 0, 0, 1, 1),
		(drawing, 5676, 5676, 0, 0, 0, 0, 1, 1),
		(drawing, 5675, 5675, 0, 0, 0, 0, 1, 1),
		(drawing, 5674, 5674, 0, 0, 0, 0, 1, 1),
		(drawing, 5673, 5673, 0, 0, 0, 0, 1, 1),
		(drawing, 5672, 5672, 0, 0, 0, 0, 1, 1),
		(drawing, 5671, 5671, 0, 0, 0, 0, 1, 1),
		(drawing, 5670, 5670, 0, 0, 0, 0, 1, 1),
		(drawing, 5669, 5669, 0, 0, 0, 0, 1, 1),
		(drawing, 5668, 5668, 0, 0, 0, 0, 1, 1),
		(drawing, 5667, 5667, 0, 0, 0, 0, 1, 1),
		(drawing, 5666, 5666, 0, 0, 0, 0, 1, 1),
		(drawing, 5665, 5665, 0, 0, 0, 0, 1, 1),
		(drawing, 5664, 5664, 0, 0, 0, 0, 1, 1),
		(drawing, 5663, 5663, 0, 0, 0, 0, 1, 1),
		(drawing, 5662, 5662, 0, 0, 0, 0, 1, 1),
		(drawing, 5661, 5661, 0, 0, 0, 0, 1, 1),
		(drawing, 5660, 5660, 0, 0, 0, 0, 1, 1),
		(drawing, 5659, 5659, 0, 0, 0, 0, 1, 1),
		(drawing, 5658, 5658, 0, 0, 0, 0, 1, 1),
		(drawing, 5657, 5657, 0, 0, 0, 0, 1, 1),
		(drawing, 5656, 5656, 0, 0, 0, 0, 1, 1),
		(drawing, 5655, 5655, 0, 0, 0, 0, 1, 1),
		(drawing, 5654, 5654, 0, 0, 0, 0, 1, 1),
		(drawing, 5653, 5653, 0, 0, 0, 0, 1, 1),
		(drawing, 5652, 5652, 0, 0, 0, 0, 1, 1),
		(drawing, 5651, 5651, 0, 0, 0, 0, 1, 1),
		(drawing, 5650, 5650, 0, 0, 0, 0, 1, 1),
		(drawing, 5649, 5649, 0, 0, 0, 0, 1, 1),
		(drawing, 5648, 5648, 0, 0, 0, 0, 1, 1),
		(drawing, 5647, 5647, 0, 0, 0, 0, 1, 1),
		(drawing, 5646, 5646, 0, 0, 0, 0, 1, 1),
		(drawing, 5645, 5645, 0, 0, 0, 0, 1, 1),
		(drawing, 5644, 5644, 0, 0, 0, 0, 1, 1),
		(drawing, 5643, 5643, 0, 0, 0, 0, 1, 1),
		(drawing, 5642, 5642, 0, 0, 0, 0, 1, 1),
		(drawing, 5641, 5641, 0, 0, 0, 0, 1, 1),
		(drawing, 5640, 5640, 0, 0, 0, 0, 1, 1),
		(drawing, 5639, 5639, 0, 0, 0, 0, 1, 1),
		(drawing, 5638, 5638, 0, 0, 0, 0, 1, 1),
		(drawing, 5637, 5637, 0, 0, 0, 0, 1, 1),
		(drawing, 5636, 5636, 0, 0, 0, 0, 1, 1),
		(drawing, 5635, 5635, 0, 0, 0, 0, 1, 1),
		(drawing, 5634, 5634, 0, 0, 0, 0, 1, 1),
		(drawing, 5633, 5633, 0, 0, 0, 0, 1, 1),
		(drawing, 5632, 5632, 0, 0, 0, 0, 1, 1),
		(drawing, 5631, 5631, 0, 0, 0, 0, 1, 1),
		(drawing, 5630, 5630, 0, 0, 0, 0, 1, 1),
		(drawing, 5629, 5629, 0, 0, 0, 0, 1, 1),
		(drawing, 5628, 5628, 0, 0, 0, 0, 1, 1),
		(drawing, 5627, 5627, 0, 0, 0, 0, 1, 1),
		(drawing, 5626, 5626, 0, 0, 0, 0, 1, 1),
		(drawing, 5625, 5625, 0, 0, 0, 0, 1, 1),
		(drawing, 5624, 5624, 0, 0, 0, 0, 1, 1),
		(drawing, 5623, 5623, 0, 0, 0, 0, 1, 1),
		(drawing, 5622, 5622, 0, 0, 0, 0, 1, 1),
		(drawing, 5621, 5621, 0, 0, 0, 0, 1, 1),
		(drawing, 5620, 5620, 0, 0, 0, 0, 1, 1),
		(drawing, 5619, 5619, 0, 0, 0, 0, 1, 1),
		(drawing, 5618, 5618, 0, 0, 0, 0, 1, 1),
		(drawing, 5617, 5617, 0, 0, 0, 0, 1, 1),
		(drawing, 5616, 5616, 0, 0, 0, 0, 1, 1),
		(drawing, 5615, 5615, 0, 0, 0, 0, 1, 1),
		(drawing, 5614, 5614, 0, 0, 0, 0, 1, 1),
		(drawing, 5613, 5613, 0, 0, 0, 0, 1, 1),
		(drawing, 5612, 5612, 0, 0, 0, 0, 1, 1),
		(drawing, 5611, 5611, 0, 0, 0, 0, 1, 1),
		(drawing, 5610, 5610, 0, 0, 0, 0, 1, 1),
		(drawing, 5609, 5609, 0, 0, 0, 0, 1, 1),
		(drawing, 5608, 5608, 0, 0, 0, 0, 1, 1),
		(drawing, 5607, 5607, 0, 0, 0, 0, 1, 1),
		(drawing, 5606, 5606, 0, 0, 0, 0, 1, 1),
		(drawing, 5605, 5605, 0, 0, 0, 0, 1, 1),
		(drawing, 5604, 5604, 0, 0, 0, 0, 1, 1),
		(drawing, 5603, 5603, 0, 0, 0, 0, 1, 1),
		(drawing, 5602, 5602, 0, 0, 0, 0, 1, 1),
		(drawing, 5601, 5601, 0, 0, 0, 0, 1, 1),
		(drawing, 5600, 5600, 0, 0, 0, 0, 1, 1),
		(drawing, 5599, 5599, 0, 0, 0, 0, 1, 1),
		(drawing, 5598, 5598, 0, 0, 0, 0, 1, 1),
		(drawing, 5597, 5597, 0, 0, 0, 0, 1, 1),
		(drawing, 5596, 5596, 0, 0, 0, 0, 1, 1),
		(drawing, 5595, 5595, 0, 0, 0, 0, 1, 1),
		(drawing, 5594, 5594, 0, 0, 0, 0, 1, 1),
		(drawing, 5593, 5593, 0, 0, 0, 0, 1, 1),
		(drawing, 5592, 5592, 0, 0, 0, 0, 1, 1),
		(drawing, 5591, 5591, 0, 0, 0, 0, 1, 1),
		(drawing, 5590, 5590, 0, 0, 0, 0, 1, 1),
		(drawing, 5589, 5589, 0, 0, 0, 0, 1, 1),
		(drawing, 5588, 5588, 0, 0, 0, 0, 1, 1),
		(drawing, 5587, 5587, 0, 0, 0, 0, 1, 1),
		(drawing, 5586, 5586, 0, 0, 0, 0, 1, 1),
		(drawing, 5585, 5585, 0, 0, 0, 0, 1, 1),
		(drawing, 5584, 5584, 0, 0, 0, 0, 1, 1),
		(drawing, 5583, 5583, 0, 0, 0, 0, 1, 1),
		(drawing, 5582, 5582, 0, 0, 0, 0, 1, 1),
		(drawing, 5581, 5581, 0, 0, 0, 0, 1, 1),
		(drawing, 5580, 5580, 0, 0, 0, 0, 1, 1),
		(drawing, 5579, 5579, 0, 0, 0, 0, 1, 1),
		(drawing, 5578, 5578, 0, 0, 0, 0, 1, 1),
		(drawing, 5577, 5577, 0, 0, 0, 0, 1, 1),
		(drawing, 5576, 5576, 0, 0, 0, 0, 1, 1),
		(drawing, 5575, 5575, 0, 0, 0, 0, 1, 1),
		(drawing, 5574, 5574, 0, 0, 0, 0, 1, 1),
		(drawing, 5573, 5573, 0, 0, 0, 0, 1, 1),
		(drawing, 5572, 5572, 0, 0, 0, 0, 1, 1),
		(drawing, 5571, 5571, 0, 0, 0, 0, 1, 1),
		(drawing, 5570, 5570, 0, 0, 0, 0, 1, 1),
		(drawing, 5569, 5569, 0, 0, 0, 0, 1, 1),
		(drawing, 5568, 5568, 0, 0, 0, 0, 1, 1),
		(drawing, 5567, 5567, 0, 0, 0, 0, 1, 1),
		(drawing, 5566, 5566, 0, 0, 0, 0, 1, 1),
		(drawing, 5565, 5565, 0, 0, 0, 0, 1, 1),
		(drawing, 5564, 5564, 0, 0, 0, 0, 1, 1),
		(drawing, 5563, 5563, 0, 0, 0, 0, 1, 1),
		(drawing, 5562, 5562, 0, 0, 0, 0, 1, 1),
		(drawing, 5561, 5561, 0, 0, 0, 0, 1, 1),
		(drawing, 5560, 5560, 0, 0, 0, 0, 1, 1),
		(drawing, 5559, 5559, 0, 0, 0, 0, 1, 1),
		(drawing, 5558, 5558, 0, 0, 0, 0, 1, 1),
		(drawing, 5557, 5557, 0, 0, 0, 0, 1, 1),
		(drawing, 5556, 5556, 0, 0, 0, 0, 1, 1),
		(drawing, 5555, 5555, 0, 0, 0, 0, 1, 1),
		(drawing, 5554, 5554, 0, 0, 0, 0, 1, 1),
		(drawing, 5553, 5553, 0, 0, 0, 0, 1, 1),
		(drawing, 5552, 5552, 0, 0, 0, 0, 1, 1),
		(drawing, 5551, 5551, 0, 0, 0, 0, 1, 1),
		(drawing, 5550, 5550, 0, 0, 0, 0, 1, 1),
		(drawing, 5549, 5549, 0, 0, 0, 0, 1, 1),
		(drawing, 5548, 5548, 0, 0, 0, 0, 1, 1),
		(drawing, 5547, 5547, 0, 0, 0, 0, 1, 1),
		(drawing, 5546, 5546, 0, 0, 0, 0, 1, 1),
		(drawing, 5545, 5545, 0, 0, 0, 0, 1, 1),
		(drawing, 5544, 5544, 0, 0, 0, 0, 1, 1),
		(drawing, 5543, 5543, 0, 0, 0, 0, 1, 1),
		(drawing, 5542, 5542, 0, 0, 0, 0, 1, 1),
		(drawing, 5541, 5541, 0, 0, 0, 0, 1, 1),
		(drawing, 5540, 5540, 0, 0, 0, 0, 1, 1),
		(drawing, 5539, 5539, 0, 0, 0, 0, 1, 1),
		(drawing, 5538, 5538, 0, 0, 0, 0, 1, 1),
		(drawing, 5537, 5537, 0, 0, 0, 0, 1, 1),
		(drawing, 5536, 5536, 0, 0, 0, 0, 1, 1),
		(drawing, 5535, 5535, 0, 0, 0, 0, 1, 1),
		(drawing, 5534, 5534, 0, 0, 0, 0, 1, 1),
		(drawing, 5533, 5533, 0, 0, 0, 0, 1, 1),
		(drawing, 5532, 5532, 0, 0, 0, 0, 1, 1),
		(drawing, 5531, 5531, 0, 0, 0, 0, 1, 1),
		(drawing, 5530, 5530, 0, 0, 0, 0, 1, 1),
		(drawing, 5529, 5529, 0, 0, 0, 0, 1, 1),
		(drawing, 5528, 5528, 0, 0, 0, 0, 1, 1),
		(drawing, 5527, 5527, 0, 0, 0, 0, 1, 1),
		(drawing, 5526, 5526, 0, 0, 0, 0, 1, 1),
		(drawing, 5525, 5525, 0, 0, 0, 0, 1, 1),
		(drawing, 5524, 5524, 0, 0, 0, 0, 1, 1),
		(drawing, 5523, 5523, 0, 0, 0, 0, 1, 1),
		(drawing, 5522, 5522, 0, 0, 0, 0, 1, 1),
		(drawing, 5521, 5521, 0, 0, 0, 0, 1, 1),
		(drawing, 5520, 5520, 0, 0, 0, 0, 1, 1),
		(drawing, 5519, 5519, 0, 0, 0, 0, 1, 1),
		(drawing, 5518, 5518, 0, 0, 0, 0, 1, 1),
		(drawing, 5517, 5517, 0, 0, 0, 0, 1, 1),
		(drawing, 5516, 5516, 0, 0, 0, 0, 1, 1),
		(drawing, 5515, 5515, 0, 0, 0, 0, 1, 1),
		(drawing, 5514, 5514, 0, 0, 0, 0, 1, 1),
		(drawing, 5513, 5513, 0, 0, 0, 0, 1, 1),
		(drawing, 5512, 5512, 0, 0, 0, 0, 1, 1),
		(drawing, 5511, 5511, 0, 0, 0, 0, 1, 1),
		(drawing, 5510, 5510, 0, 0, 0, 0, 1, 1),
		(drawing, 5509, 5509, 0, 0, 0, 0, 1, 1),
		(drawing, 5508, 5508, 0, 0, 0, 0, 1, 1),
		(drawing, 5507, 5507, 0, 0, 0, 0, 1, 1),
		(drawing, 5506, 5506, 0, 0, 0, 0, 1, 1),
		(drawing, 5505, 5505, 0, 0, 0, 0, 1, 1),
		(drawing, 5504, 5504, 0, 0, 0, 0, 1, 1),
		(drawing, 5503, 5503, 0, 0, 0, 0, 1, 1),
		(drawing, 5502, 5502, 0, 0, 0, 0, 1, 1),
		(drawing, 5501, 5501, 0, 0, 0, 0, 1, 1),
		(drawing, 5500, 5500, 0, 0, 0, 0, 1, 1),
		(drawing, 5499, 5499, 0, 0, 0, 0, 1, 1),
		(drawing, 5498, 5498, 0, 0, 0, 0, 1, 1),
		(drawing, 5497, 5497, 0, 0, 0, 0, 1, 1),
		(drawing, 5496, 5496, 0, 0, 0, 0, 1, 1),
		(drawing, 5495, 5495, 0, 0, 0, 0, 1, 1),
		(drawing, 5494, 5494, 0, 0, 0, 0, 1, 1),
		(drawing, 5493, 5493, 0, 0, 0, 0, 1, 1),
		(drawing, 5492, 5492, 0, 0, 0, 0, 1, 1),
		(drawing, 5491, 5491, 0, 0, 0, 0, 1, 1),
		(drawing, 5490, 5490, 0, 0, 0, 0, 1, 1),
		(drawing, 5489, 5489, 0, 0, 0, 0, 1, 1),
		(drawing, 5488, 5488, 0, 0, 0, 0, 1, 1),
		(drawing, 5487, 5487, 0, 0, 0, 0, 1, 1),
		(drawing, 5486, 5486, 0, 0, 0, 0, 1, 1),
		(drawing, 5485, 5485, 0, 0, 0, 0, 1, 1),
		(drawing, 5484, 5484, 0, 0, 0, 0, 1, 1),
		(drawing, 5483, 5483, 0, 0, 0, 0, 1, 1),
		(drawing, 5482, 5482, 0, 0, 0, 0, 1, 1),
		(drawing, 5481, 5481, 0, 0, 0, 0, 1, 1),
		(drawing, 5480, 5480, 0, 0, 0, 0, 1, 1),
		(drawing, 5479, 5479, 0, 0, 0, 0, 1, 1),
		(drawing, 5478, 5478, 0, 0, 0, 0, 1, 1),
		(drawing, 5477, 5477, 0, 0, 0, 0, 1, 1),
		(drawing, 5476, 5476, 0, 0, 0, 0, 1, 1),
		(drawing, 5475, 5475, 0, 0, 0, 0, 1, 1),
		(drawing, 5474, 5474, 0, 0, 0, 0, 1, 1),
		(drawing, 5473, 5473, 0, 0, 0, 0, 1, 1),
		(drawing, 5472, 5472, 0, 0, 0, 0, 1, 1),
		(drawing, 5471, 5471, 0, 0, 0, 0, 1, 1),
		(drawing, 5470, 5470, 0, 0, 0, 0, 1, 1),
		(drawing, 5469, 5469, 0, 0, 0, 0, 1, 1),
		(drawing, 5468, 5468, 0, 0, 0, 0, 1, 1),
		(drawing, 5467, 5467, 0, 0, 0, 0, 1, 1),
		(drawing, 5466, 5466, 0, 0, 0, 0, 1, 1),
		(drawing, 5465, 5465, 0, 0, 0, 0, 1, 1),
		(drawing, 5464, 5464, 0, 0, 0, 0, 1, 1),
		(drawing, 5463, 5463, 0, 0, 0, 0, 1, 1),
		(drawing, 5462, 5462, 0, 0, 0, 0, 1, 1),
		(drawing, 5461, 5461, 0, 0, 0, 0, 1, 1),
		(drawing, 5460, 5460, 0, 0, 0, 0, 1, 1),
		(drawing, 5459, 5459, 0, 0, 0, 0, 1, 1),
		(drawing, 5458, 5458, 0, 0, 0, 0, 1, 1),
		(drawing, 5457, 5457, 0, 0, 0, 0, 1, 1),
		(drawing, 5456, 5456, 0, 0, 0, 0, 1, 1),
		(drawing, 5455, 5455, 0, 0, 0, 0, 1, 1),
		(drawing, 5454, 5454, 0, 0, 0, 0, 1, 1),
		(drawing, 5453, 5453, 0, 0, 0, 0, 1, 1),
		(drawing, 5452, 5452, 0, 0, 0, 0, 1, 1),
		(drawing, 5451, 5451, 0, 0, 0, 0, 1, 1),
		(drawing, 5450, 5450, 0, 0, 0, 0, 1, 1),
		(drawing, 5449, 5449, 0, 0, 0, 0, 1, 1),
		(drawing, 5448, 5448, 0, 0, 0, 0, 1, 1),
		(drawing, 5447, 5447, 0, 0, 0, 0, 1, 1),
		(drawing, 5446, 5446, 0, 0, 0, 0, 1, 1),
		(drawing, 5445, 5445, 0, 0, 0, 0, 1, 1),
		(drawing, 5444, 5444, 0, 0, 0, 0, 1, 1),
		(drawing, 5443, 5443, 0, 0, 0, 0, 1, 1),
		(drawing, 5442, 5442, 0, 0, 0, 0, 1, 1),
		(drawing, 5441, 5441, 0, 0, 0, 0, 1, 1),
		(drawing, 5440, 5440, 0, 0, 0, 0, 1, 1),
		(drawing, 5439, 5439, 0, 0, 0, 0, 1, 1),
		(drawing, 5438, 5438, 0, 0, 0, 0, 1, 1),
		(drawing, 5437, 5437, 0, 0, 0, 0, 1, 1),
		(drawing, 5436, 5436, 0, 0, 0, 0, 1, 1),
		(drawing, 5435, 5435, 0, 0, 0, 0, 1, 1),
		(drawing, 5434, 5434, 0, 0, 0, 0, 1, 1),
		(drawing, 5433, 5433, 0, 0, 0, 0, 1, 1),
		(drawing, 5432, 5432, 0, 0, 0, 0, 1, 1),
		(drawing, 5431, 5431, 0, 0, 0, 0, 1, 1),
		(drawing, 5430, 5430, 0, 0, 0, 0, 1, 1),
		(drawing, 5429, 5429, 0, 0, 0, 0, 1, 1),
		(drawing, 5428, 5428, 0, 0, 0, 0, 1, 1),
		(drawing, 5427, 5427, 0, 0, 0, 0, 1, 1),
		(drawing, 5426, 5426, 0, 0, 0, 0, 1, 1),
		(drawing, 5425, 5425, 0, 0, 0, 0, 1, 1),
		(drawing, 5424, 5424, 0, 0, 0, 0, 1, 1),
		(drawing, 5423, 5423, 0, 0, 0, 0, 1, 1),
		(drawing, 5422, 5422, 0, 0, 0, 0, 1, 1),
		(drawing, 5421, 5421, 0, 0, 0, 0, 1, 1),
		(drawing, 5420, 5420, 0, 0, 0, 0, 1, 1),
		(drawing, 5419, 5419, 0, 0, 0, 0, 1, 1),
		(drawing, 5418, 5418, 0, 0, 0, 0, 1, 1),
		(drawing, 5417, 5417, 0, 0, 0, 0, 1, 1),
		(drawing, 5416, 5416, 0, 0, 0, 0, 1, 1),
		(drawing, 5415, 5415, 0, 0, 0, 0, 1, 1),
		(drawing, 5414, 5414, 0, 0, 0, 0, 1, 1),
		(drawing, 5413, 5413, 0, 0, 0, 0, 1, 1),
		(drawing, 5412, 5412, 0, 0, 0, 0, 1, 1),
		(drawing, 5411, 5411, 0, 0, 0, 0, 1, 1),
		(drawing, 5410, 5410, 0, 0, 0, 0, 1, 1),
		(drawing, 5409, 5409, 0, 0, 0, 0, 1, 1),
		(drawing, 5408, 5408, 0, 0, 0, 0, 1, 1),
		(drawing, 5407, 5407, 0, 0, 0, 0, 1, 1),
		(drawing, 5406, 5406, 0, 0, 0, 0, 1, 1),
		(drawing, 5405, 5405, 0, 0, 0, 0, 1, 1),
		(drawing, 5404, 5404, 0, 0, 0, 0, 1, 1),
		(drawing, 5403, 5403, 0, 0, 0, 0, 1, 1),
		(drawing, 5402, 5402, 0, 0, 0, 0, 1, 1),
		(drawing, 5401, 5401, 0, 0, 0, 0, 1, 1),
		(drawing, 5400, 5400, 0, 0, 0, 0, 1, 1),
		(drawing, 5399, 5399, 0, 0, 0, 0, 1, 1),
		(drawing, 5398, 5398, 0, 0, 0, 0, 1, 1),
		(drawing, 5397, 5397, 0, 0, 0, 0, 1, 1),
		(drawing, 5396, 5396, 0, 0, 0, 0, 1, 1),
		(drawing, 5395, 5395, 0, 0, 0, 0, 1, 1),
		(drawing, 5394, 5394, 0, 0, 0, 0, 1, 1),
		(drawing, 5393, 5393, 0, 0, 0, 0, 1, 1),
		(drawing, 5392, 5392, 0, 0, 0, 0, 1, 1),
		(drawing, 5391, 5391, 0, 0, 0, 0, 1, 1),
		(drawing, 5390, 5390, 0, 0, 0, 0, 1, 1),
		(drawing, 5389, 5389, 0, 0, 0, 0, 1, 1),
		(drawing, 5388, 5388, 0, 0, 0, 0, 1, 1),
		(drawing, 5387, 5387, 0, 0, 0, 0, 1, 1),
		(drawing, 5386, 5386, 0, 0, 0, 0, 1, 1),
		(drawing, 5385, 5385, 0, 0, 0, 0, 1, 1),
		(drawing, 5384, 5384, 0, 0, 0, 0, 1, 1),
		(drawing, 5383, 5383, 0, 0, 0, 0, 1, 1),
		(drawing, 5382, 5382, 0, 0, 0, 0, 1, 1),
		(drawing, 5381, 5381, 0, 0, 0, 0, 1, 1),
		(drawing, 5380, 5380, 0, 0, 0, 0, 1, 1),
		(drawing, 5379, 5379, 0, 0, 0, 0, 1, 1),
		(drawing, 5378, 5378, 0, 0, 0, 0, 1, 1),
		(drawing, 5377, 5377, 0, 0, 0, 0, 1, 1),
		(drawing, 5376, 5376, 0, 0, 0, 0, 1, 1),
		(drawing, 5375, 5375, 0, 0, 0, 0, 1, 1),
		(drawing, 5374, 5374, 0, 0, 0, 0, 1, 1),
		(drawing, 5373, 5373, 0, 0, 0, 0, 1, 1),
		(drawing, 5372, 5372, 0, 0, 0, 0, 1, 1),
		(drawing, 5371, 5371, 0, 0, 0, 0, 1, 1),
		(drawing, 5370, 5370, 0, 0, 0, 0, 1, 1),
		(drawing, 5369, 5369, 0, 0, 0, 0, 1, 1),
		(drawing, 5368, 5368, 0, 0, 0, 0, 1, 1),
		(drawing, 5367, 5367, 0, 0, 0, 0, 1, 1),
		(drawing, 5366, 5366, 0, 0, 0, 0, 1, 1),
		(drawing, 5365, 5365, 0, 0, 0, 0, 1, 1),
		(drawing, 5364, 5364, 0, 0, 0, 0, 1, 1),
		(drawing, 5363, 5363, 0, 0, 0, 0, 1, 1),
		(drawing, 5362, 5362, 0, 0, 0, 0, 1, 1),
		(drawing, 5361, 5361, 0, 0, 0, 0, 1, 1),
		(drawing, 5360, 5360, 0, 0, 0, 0, 1, 1),
		(drawing, 5359, 5359, 0, 0, 0, 0, 1, 1),
		(drawing, 5358, 5358, 0, 0, 0, 0, 1, 1),
		(drawing, 5357, 5357, 0, 0, 0, 0, 1, 1),
		(drawing, 5356, 5356, 0, 0, 0, 0, 1, 1),
		(drawing, 5355, 5355, 0, 0, 0, 0, 1, 1),
		(drawing, 5354, 5354, 0, 0, 0, 0, 1, 1),
		(drawing, 5353, 5353, 0, 0, 0, 0, 1, 1),
		(drawing, 5352, 5352, 0, 0, 0, 0, 1, 1),
		(drawing, 5351, 5351, 0, 0, 0, 0, 1, 1),
		(drawing, 5350, 5350, 0, 0, 0, 0, 1, 1),
		(drawing, 5349, 5349, 0, 0, 0, 0, 1, 1),
		(drawing, 5348, 5348, 0, 0, 0, 0, 1, 1),
		(drawing, 5347, 5347, 0, 0, 0, 0, 1, 1),
		(drawing, 5346, 5346, 0, 0, 0, 0, 1, 1),
		(drawing, 5345, 5345, 0, 0, 0, 0, 1, 1),
		(drawing, 5344, 5344, 0, 0, 0, 0, 1, 1),
		(drawing, 5343, 5343, 0, 0, 0, 0, 1, 1),
		(drawing, 5342, 5342, 0, 0, 0, 0, 1, 1),
		(drawing, 5341, 5341, 0, 0, 0, 0, 1, 1),
		(drawing, 5340, 5340, 0, 0, 0, 0, 1, 1),
		(drawing, 5339, 5339, 0, 0, 0, 0, 1, 1),
		(drawing, 5338, 5338, 0, 0, 0, 0, 1, 1),
		(drawing, 5337, 5337, 0, 0, 0, 0, 1, 1),
		(drawing, 5336, 5336, 0, 0, 0, 0, 1, 1),
		(drawing, 5335, 5335, 0, 0, 0, 0, 1, 1),
		(drawing, 5334, 5334, 0, 0, 0, 0, 1, 1),
		(drawing, 5333, 5333, 0, 0, 0, 0, 1, 1),
		(drawing, 5332, 5332, 0, 0, 0, 0, 1, 1),
		(drawing, 5331, 5331, 0, 0, 0, 0, 1, 1),
		(drawing, 5330, 5330, 0, 0, 0, 0, 1, 1),
		(drawing, 5329, 5329, 0, 0, 0, 0, 1, 1),
		(drawing, 5328, 5328, 0, 0, 0, 0, 1, 1),
		(drawing, 5327, 5327, 0, 0, 0, 0, 1, 1),
		(drawing, 5326, 5326, 0, 0, 0, 0, 1, 1),
		(drawing, 5325, 5325, 0, 0, 0, 0, 1, 1),
		(drawing, 5324, 5324, 0, 0, 0, 0, 1, 1),
		(drawing, 5323, 5323, 0, 0, 0, 0, 1, 1),
		(drawing, 5322, 5322, 0, 0, 0, 0, 1, 1),
		(drawing, 5321, 5321, 0, 0, 0, 0, 1, 1),
		(drawing, 5320, 5320, 0, 0, 0, 0, 1, 1),
		(drawing, 5319, 5319, 0, 0, 0, 0, 1, 1),
		(drawing, 5318, 5318, 0, 0, 0, 0, 1, 1),
		(drawing, 5317, 5317, 0, 0, 0, 0, 1, 1),
		(drawing, 5316, 5316, 0, 0, 0, 0, 1, 1),
		(drawing, 5315, 5315, 0, 0, 0, 0, 1, 1),
		(drawing, 5314, 5314, 0, 0, 0, 0, 1, 1),
		(drawing, 5313, 5313, 0, 0, 0, 0, 1, 1),
		(drawing, 5312, 5312, 0, 0, 0, 0, 1, 1),
		(drawing, 5311, 5311, 0, 0, 0, 0, 1, 1),
		(drawing, 5310, 5310, 0, 0, 0, 0, 1, 1),
		(drawing, 5309, 5309, 0, 0, 0, 0, 1, 1),
		(drawing, 5308, 5308, 0, 0, 0, 0, 1, 1),
		(drawing, 5307, 5307, 0, 0, 0, 0, 1, 1),
		(drawing, 5306, 5306, 0, 0, 0, 0, 1, 1),
		(drawing, 5305, 5305, 0, 0, 0, 0, 1, 1),
		(drawing, 5304, 5304, 0, 0, 0, 0, 1, 1),
		(drawing, 5303, 5303, 0, 0, 0, 0, 1, 1),
		(drawing, 5302, 5302, 0, 0, 0, 0, 1, 1),
		(drawing, 5301, 5301, 0, 0, 0, 0, 1, 1),
		(drawing, 5300, 5300, 0, 0, 0, 0, 1, 1),
		(drawing, 5299, 5299, 0, 0, 0, 0, 1, 1),
		(drawing, 5298, 5298, 0, 0, 0, 0, 1, 1),
		(drawing, 5297, 5297, 0, 0, 0, 0, 1, 1),
		(drawing, 5296, 5296, 0, 0, 0, 0, 1, 1),
		(drawing, 5295, 5295, 0, 0, 0, 0, 1, 1),
		(drawing, 5294, 5294, 0, 0, 0, 0, 1, 1),
		(drawing, 5293, 5293, 0, 0, 0, 0, 1, 1),
		(drawing, 5292, 5292, 0, 0, 0, 0, 1, 1),
		(drawing, 5291, 5291, 0, 0, 0, 0, 1, 1),
		(drawing, 5290, 5290, 0, 0, 0, 0, 1, 1),
		(drawing, 5289, 5289, 0, 0, 0, 0, 1, 1),
		(drawing, 5288, 5288, 0, 0, 0, 0, 1, 1),
		(drawing, 5287, 5287, 0, 0, 0, 0, 1, 1),
		(drawing, 5286, 5286, 0, 0, 0, 0, 1, 1),
		(drawing, 5285, 5285, 0, 0, 0, 0, 1, 1),
		(drawing, 5284, 5284, 0, 0, 0, 0, 1, 1),
		(drawing, 5283, 5283, 0, 0, 0, 0, 1, 1),
		(drawing, 5282, 5282, 0, 0, 0, 0, 1, 1),
		(drawing, 5281, 5281, 0, 0, 0, 0, 1, 1),
		(drawing, 5280, 5280, 0, 0, 0, 0, 1, 1),
		(drawing, 5279, 5279, 0, 0, 0, 0, 1, 1),
		(drawing, 5278, 5278, 0, 0, 0, 0, 1, 1),
		(drawing, 5277, 5277, 0, 0, 0, 0, 1, 1),
		(drawing, 5276, 5276, 0, 0, 0, 0, 1, 1),
		(drawing, 5275, 5275, 0, 0, 0, 0, 1, 1),
		(drawing, 5274, 5274, 0, 0, 0, 0, 1, 1),
		(drawing, 5273, 5273, 0, 0, 0, 0, 1, 1),
		(drawing, 5272, 5272, 0, 0, 0, 0, 1, 1),
		(drawing, 5271, 5271, 0, 0, 0, 0, 1, 1),
		(drawing, 5270, 5270, 0, 0, 0, 0, 1, 1),
		(drawing, 5269, 5269, 0, 0, 0, 0, 1, 1),
		(drawing, 5268, 5268, 0, 0, 0, 0, 1, 1),
		(drawing, 5267, 5267, 0, 0, 0, 0, 1, 1),
		(drawing, 5266, 5266, 0, 0, 0, 0, 1, 1),
		(drawing, 5265, 5265, 0, 0, 0, 0, 1, 1),
		(drawing, 5264, 5264, 0, 0, 0, 0, 1, 1),
		(drawing, 5263, 5263, 0, 0, 0, 0, 1, 1),
		(drawing, 5262, 5262, 0, 0, 0, 0, 1, 1),
		(drawing, 5261, 5261, 0, 0, 0, 0, 1, 1),
		(drawing, 5260, 5260, 0, 0, 0, 0, 1, 1),
		(drawing, 5259, 5259, 0, 0, 0, 0, 1, 1),
		(drawing, 5258, 5258, 0, 0, 0, 0, 1, 1),
		(drawing, 5257, 5257, 0, 0, 0, 0, 1, 1),
		(drawing, 5256, 5256, 0, 0, 0, 0, 1, 1),
		(drawing, 5255, 5255, 0, 0, 0, 0, 1, 1),
		(drawing, 5254, 5254, 0, 0, 0, 0, 1, 1),
		(drawing, 5253, 5253, 0, 0, 0, 0, 1, 1),
		(drawing, 5252, 5252, 0, 0, 0, 0, 1, 1),
		(drawing, 5251, 5251, 0, 0, 0, 0, 1, 1),
		(drawing, 5250, 5250, 0, 0, 0, 0, 1, 1),
		(drawing, 5249, 5249, 0, 0, 0, 0, 1, 1),
		(drawing, 5248, 5248, 0, 0, 0, 0, 1, 1),
		(drawing, 5247, 5247, 0, 0, 0, 0, 1, 1),
		(drawing, 5246, 5246, 0, 0, 0, 0, 1, 1),
		(drawing, 5245, 5245, 0, 0, 0, 0, 1, 1),
		(drawing, 5244, 5244, 0, 0, 0, 0, 1, 1),
		(drawing, 5243, 5243, 0, 0, 0, 0, 1, 1),
		(drawing, 5242, 5242, 0, 0, 0, 0, 1, 1),
		(drawing, 5241, 5241, 0, 0, 0, 0, 1, 1),
		(drawing, 5240, 5240, 0, 0, 0, 0, 1, 1),
		(drawing, 5239, 5239, 0, 0, 0, 0, 1, 1),
		(drawing, 5238, 5238, 0, 0, 0, 0, 1, 1),
		(drawing, 5237, 5237, 0, 0, 0, 0, 1, 1),
		(drawing, 5236, 5236, 0, 0, 0, 0, 1, 1),
		(drawing, 5235, 5235, 0, 0, 0, 0, 1, 1),
		(drawing, 5234, 5234, 0, 0, 0, 0, 1, 1),
		(drawing, 5233, 5233, 0, 0, 0, 0, 1, 1),
		(drawing, 5232, 5232, 0, 0, 0, 0, 1, 1),
		(drawing, 5231, 5231, 0, 0, 0, 0, 1, 1),
		(drawing, 5230, 5230, 0, 0, 0, 0, 1, 1),
		(drawing, 5229, 5229, 0, 0, 0, 0, 1, 1),
		(drawing, 5228, 5228, 0, 0, 0, 0, 1, 1),
		(drawing, 5227, 5227, 0, 0, 0, 0, 1, 1),
		(drawing, 5226, 5226, 0, 0, 0, 0, 1, 1),
		(drawing, 5225, 5225, 0, 0, 0, 0, 1, 1),
		(drawing, 5224, 5224, 0, 0, 0, 0, 1, 1),
		(drawing, 5223, 5223, 0, 0, 0, 0, 1, 1),
		(drawing, 5222, 5222, 0, 0, 0, 0, 1, 1),
		(drawing, 5221, 5221, 0, 0, 0, 0, 1, 1),
		(drawing, 5220, 5220, 0, 0, 0, 0, 1, 1),
		(drawing, 5219, 5219, 0, 0, 0, 0, 1, 1),
		(drawing, 5218, 5218, 0, 0, 0, 0, 1, 1),
		(drawing, 5217, 5217, 0, 0, 0, 0, 1, 1),
		(drawing, 5216, 5216, 0, 0, 0, 0, 1, 1),
		(drawing, 5215, 5215, 0, 0, 0, 0, 1, 1),
		(drawing, 5214, 5214, 0, 0, 0, 0, 1, 1),
		(drawing, 5213, 5213, 0, 0, 0, 0, 1, 1),
		(drawing, 5212, 5212, 0, 0, 0, 0, 1, 1),
		(drawing, 5211, 5211, 0, 0, 0, 0, 1, 1),
		(drawing, 5210, 5210, 0, 0, 0, 0, 1, 1),
		(drawing, 5209, 5209, 0, 0, 0, 0, 1, 1),
		(drawing, 5208, 5208, 0, 0, 0, 0, 1, 1),
		(drawing, 5207, 5207, 0, 0, 0, 0, 1, 1),
		(drawing, 5206, 5206, 0, 0, 0, 0, 1, 1),
		(drawing, 5205, 5205, 0, 0, 0, 0, 1, 1),
		(drawing, 5204, 5204, 0, 0, 0, 0, 1, 1),
		(drawing, 5203, 5203, 0, 0, 0, 0, 1, 1),
		(drawing, 5202, 5202, 0, 0, 0, 0, 1, 1),
		(drawing, 5201, 5201, 0, 0, 0, 0, 1, 1),
		(drawing, 5200, 5200, 0, 0, 0, 0, 1, 1),
		(drawing, 5199, 5199, 0, 0, 0, 0, 1, 1),
		(drawing, 5198, 5198, 0, 0, 0, 0, 1, 1),
		(drawing, 5197, 5197, 0, 0, 0, 0, 1, 1),
		(drawing, 5196, 5196, 0, 0, 0, 0, 1, 1),
		(drawing, 5195, 5195, 0, 0, 0, 0, 1, 1),
		(drawing, 5194, 5194, 0, 0, 0, 0, 1, 1),
		(drawing, 5193, 5193, 0, 0, 0, 0, 1, 1),
		(drawing, 5192, 5192, 0, 0, 0, 0, 1, 1),
		(drawing, 5191, 5191, 0, 0, 0, 0, 1, 1),
		(drawing, 5190, 5190, 0, 0, 0, 0, 1, 1),
		(drawing, 5189, 5189, 0, 0, 0, 0, 1, 1),
		(drawing, 5188, 5188, 0, 0, 0, 0, 1, 1),
		(drawing, 5187, 5187, 0, 0, 0, 0, 1, 1),
		(drawing, 5186, 5186, 0, 0, 0, 0, 1, 1),
		(drawing, 5185, 5185, 0, 0, 0, 0, 1, 1),
		(drawing, 5184, 5184, 0, 0, 0, 0, 1, 1),
		(drawing, 5183, 5183, 0, 0, 0, 0, 1, 1),
		(drawing, 5182, 5182, 0, 0, 0, 0, 1, 1),
		(drawing, 5181, 5181, 0, 0, 0, 0, 1, 1),
		(drawing, 5180, 5180, 0, 0, 0, 0, 1, 1),
		(drawing, 5179, 5179, 0, 0, 0, 0, 1, 1),
		(drawing, 5178, 5178, 0, 0, 0, 0, 1, 1),
		(drawing, 5177, 5177, 0, 0, 0, 0, 1, 1),
		(drawing, 5176, 5176, 0, 0, 0, 0, 1, 1),
		(drawing, 5175, 5175, 0, 0, 0, 0, 1, 1),
		(drawing, 5174, 5174, 0, 0, 0, 0, 1, 1),
		(drawing, 5173, 5173, 0, 0, 0, 0, 1, 1),
		(drawing, 5172, 5172, 0, 0, 0, 0, 1, 1),
		(drawing, 5171, 5171, 0, 0, 0, 0, 1, 1),
		(drawing, 5170, 5170, 0, 0, 0, 0, 1, 1),
		(drawing, 5169, 5169, 0, 0, 0, 0, 1, 1),
		(drawing, 5168, 5168, 0, 0, 0, 0, 1, 1),
		(drawing, 5167, 5167, 0, 0, 0, 0, 1, 1),
		(drawing, 5166, 5166, 0, 0, 0, 0, 1, 1),
		(drawing, 5165, 5165, 0, 0, 0, 0, 1, 1),
		(drawing, 5164, 5164, 0, 0, 0, 0, 1, 1),
		(drawing, 5163, 5163, 0, 0, 0, 0, 1, 1),
		(drawing, 5162, 5162, 0, 0, 0, 0, 1, 1),
		(drawing, 5161, 5161, 0, 0, 0, 0, 1, 1),
		(drawing, 5160, 5160, 0, 0, 0, 0, 1, 1),
		(drawing, 5159, 5159, 0, 0, 0, 0, 1, 1),
		(drawing, 5158, 5158, 0, 0, 0, 0, 1, 1),
		(drawing, 5157, 5157, 0, 0, 0, 0, 1, 1),
		(drawing, 5156, 5156, 0, 0, 0, 0, 1, 1),
		(drawing, 5155, 5155, 0, 0, 0, 0, 1, 1),
		(drawing, 5154, 5154, 0, 0, 0, 0, 1, 1),
		(drawing, 5153, 5153, 0, 0, 0, 0, 1, 1),
		(drawing, 5152, 5152, 0, 0, 0, 0, 1, 1),
		(drawing, 5151, 5151, 0, 0, 0, 0, 1, 1),
		(drawing, 5150, 5150, 0, 0, 0, 0, 1, 1),
		(drawing, 5149, 5149, 0, 0, 0, 0, 1, 1),
		(drawing, 5148, 5148, 0, 0, 0, 0, 1, 1),
		(drawing, 5147, 5147, 0, 0, 0, 0, 1, 1),
		(drawing, 5146, 5146, 0, 0, 0, 0, 1, 1),
		(drawing, 5145, 5145, 0, 0, 0, 0, 1, 1),
		(drawing, 5144, 5144, 0, 0, 0, 0, 1, 1),
		(drawing, 5143, 5143, 0, 0, 0, 0, 1, 1),
		(drawing, 5142, 5142, 0, 0, 0, 0, 1, 1),
		(drawing, 5141, 5141, 0, 0, 0, 0, 1, 1),
		(drawing, 5140, 5140, 0, 0, 0, 0, 1, 1),
		(drawing, 5139, 5139, 0, 0, 0, 0, 1, 1),
		(drawing, 5138, 5138, 0, 0, 0, 0, 1, 1),
		(drawing, 5137, 5137, 0, 0, 0, 0, 1, 1),
		(drawing, 5136, 5136, 0, 0, 0, 0, 1, 1),
		(drawing, 5135, 5135, 0, 0, 0, 0, 1, 1),
		(drawing, 5134, 5134, 0, 0, 0, 0, 1, 1),
		(drawing, 5133, 5133, 0, 0, 0, 0, 1, 1),
		(drawing, 5132, 5132, 0, 0, 0, 0, 1, 1),
		(drawing, 5131, 5131, 0, 0, 0, 0, 1, 1),
		(drawing, 5130, 5130, 0, 0, 0, 0, 1, 1),
		(drawing, 5129, 5129, 0, 0, 0, 0, 1, 1),
		(drawing, 5128, 5128, 0, 0, 0, 0, 1, 1),
		(drawing, 5127, 5127, 0, 0, 0, 0, 1, 1),
		(drawing, 5126, 5126, 0, 0, 0, 0, 1, 1),
		(drawing, 5125, 5125, 0, 0, 0, 0, 1, 1),
		(drawing, 5124, 5124, 0, 0, 0, 0, 1, 1),
		(drawing, 5123, 5123, 0, 0, 0, 0, 1, 1),
		(drawing, 5122, 5122, 0, 0, 0, 0, 1, 1),
		(drawing, 5121, 5121, 0, 0, 0, 0, 1, 1),
		(drawing, 5120, 5120, 0, 0, 0, 0, 1, 1),
		(drawing, 5119, 5119, 0, 0, 0, 0, 1, 1),
		(drawing, 5118, 5118, 0, 0, 0, 0, 1, 1),
		(drawing, 5117, 5117, 0, 0, 0, 0, 1, 1),
		(drawing, 5116, 5116, 0, 0, 0, 0, 1, 1),
		(drawing, 5115, 5115, 0, 0, 0, 0, 1, 1),
		(drawing, 5114, 5114, 0, 0, 0, 0, 1, 1),
		(drawing, 5113, 5113, 0, 0, 0, 0, 1, 1),
		(drawing, 5112, 5112, 0, 0, 0, 0, 1, 1),
		(drawing, 5111, 5111, 0, 0, 0, 0, 1, 1),
		(drawing, 5110, 5110, 0, 0, 0, 0, 1, 1),
		(drawing, 5109, 5109, 0, 0, 0, 0, 1, 1),
		(drawing, 5108, 5108, 0, 0, 0, 0, 1, 1),
		(drawing, 5107, 5107, 0, 0, 0, 0, 1, 1),
		(drawing, 5106, 5106, 0, 0, 0, 0, 1, 1),
		(drawing, 5105, 5105, 0, 0, 0, 0, 1, 1),
		(drawing, 5104, 5104, 0, 0, 0, 0, 1, 1),
		(drawing, 5103, 5103, 0, 0, 0, 0, 1, 1),
		(drawing, 5102, 5102, 0, 0, 0, 0, 1, 1),
		(drawing, 5101, 5101, 0, 0, 0, 0, 1, 1),
		(drawing, 5100, 5100, 0, 0, 0, 0, 1, 1),
		(drawing, 5099, 5099, 0, 0, 0, 0, 1, 1),
		(drawing, 5098, 5098, 0, 0, 0, 0, 1, 1),
		(drawing, 5097, 5097, 0, 0, 0, 0, 1, 1),
		(drawing, 5096, 5096, 0, 0, 0, 0, 1, 1),
		(drawing, 5095, 5095, 0, 0, 0, 0, 1, 1),
		(drawing, 5094, 5094, 0, 0, 0, 0, 1, 1),
		(drawing, 5093, 5093, 0, 0, 0, 0, 1, 1),
		(drawing, 5092, 5092, 0, 0, 0, 0, 1, 1),
		(drawing, 5091, 5091, 0, 0, 0, 0, 1, 1),
		(drawing, 5090, 5090, 0, 0, 0, 0, 1, 1),
		(drawing, 5089, 5089, 0, 0, 0, 0, 1, 1),
		(drawing, 5088, 5088, 0, 0, 0, 0, 1, 1),
		(drawing, 5087, 5087, 0, 0, 0, 0, 1, 1),
		(drawing, 5086, 5086, 0, 0, 0, 0, 1, 1),
		(drawing, 5085, 5085, 0, 0, 0, 0, 1, 1),
		(drawing, 5084, 5084, 0, 0, 0, 0, 1, 1),
		(drawing, 5083, 5083, 0, 0, 0, 0, 1, 1),
		(drawing, 5082, 5082, 0, 0, 0, 0, 1, 1),
		(drawing, 5081, 5081, 0, 0, 0, 0, 1, 1),
		(drawing, 5080, 5080, 0, 0, 0, 0, 1, 1),
		(drawing, 5079, 5079, 0, 0, 0, 0, 1, 1),
		(drawing, 5078, 5078, 0, 0, 0, 0, 1, 1),
		(drawing, 5077, 5077, 0, 0, 0, 0, 1, 1),
		(drawing, 5076, 5076, 0, 0, 0, 0, 1, 1),
		(drawing, 5075, 5075, 0, 0, 0, 0, 1, 1),
		(drawing, 5074, 5074, 0, 0, 0, 0, 1, 1),
		(drawing, 5073, 5073, 0, 0, 0, 0, 1, 1),
		(drawing, 5072, 5072, 0, 0, 0, 0, 1, 1),
		(drawing, 5071, 5071, 0, 0, 0, 0, 1, 1),
		(drawing, 5070, 5070, 0, 0, 0, 0, 1, 1),
		(drawing, 5069, 5069, 0, 0, 0, 0, 1, 1),
		(drawing, 5068, 5068, 0, 0, 0, 0, 1, 1),
		(drawing, 5067, 5067, 0, 0, 0, 0, 1, 1),
		(drawing, 5066, 5066, 0, 0, 0, 0, 1, 1),
		(drawing, 5065, 5065, 0, 0, 0, 0, 1, 1),
		(drawing, 5064, 5064, 0, 0, 0, 0, 1, 1),
		(drawing, 5063, 5063, 0, 0, 0, 0, 1, 1),
		(drawing, 5062, 5062, 0, 0, 0, 0, 1, 1),
		(drawing, 5061, 5061, 0, 0, 0, 0, 1, 1),
		(drawing, 5060, 5060, 0, 0, 0, 0, 1, 1),
		(drawing, 5059, 5059, 0, 0, 0, 0, 1, 1),
		(drawing, 5058, 5058, 0, 0, 0, 0, 1, 1),
		(drawing, 5057, 5057, 0, 0, 0, 0, 1, 1),
		(drawing, 5056, 5056, 0, 0, 0, 0, 1, 1),
		(drawing, 5055, 5055, 0, 0, 0, 0, 1, 1),
		(drawing, 5054, 5054, 0, 0, 0, 0, 1, 1),
		(drawing, 5053, 5053, 0, 0, 0, 0, 1, 1),
		(drawing, 5052, 5052, 0, 0, 0, 0, 1, 1),
		(drawing, 5051, 5051, 0, 0, 0, 0, 1, 1),
		(drawing, 5050, 5050, 0, 0, 0, 0, 1, 1),
		(drawing, 5049, 5049, 0, 0, 0, 0, 1, 1),
		(drawing, 5048, 5048, 0, 0, 0, 0, 1, 1),
		(drawing, 5047, 5047, 0, 0, 0, 0, 1, 1),
		(drawing, 5046, 5046, 0, 0, 0, 0, 1, 1),
		(drawing, 5045, 5045, 0, 0, 0, 0, 1, 1),
		(drawing, 5044, 5044, 0, 0, 0, 0, 1, 1),
		(drawing, 5043, 5043, 0, 0, 0, 0, 1, 1),
		(drawing, 5042, 5042, 0, 0, 0, 0, 1, 1),
		(drawing, 5041, 5041, 0, 0, 0, 0, 1, 1),
		(drawing, 5040, 5040, 0, 0, 0, 0, 1, 1),
		(drawing, 5039, 5039, 0, 0, 0, 0, 1, 1),
		(drawing, 5038, 5038, 0, 0, 0, 0, 1, 1),
		(drawing, 5037, 5037, 0, 0, 0, 0, 1, 1),
		(drawing, 5036, 5036, 0, 0, 0, 0, 1, 1),
		(drawing, 5035, 5035, 0, 0, 0, 0, 1, 1),
		(drawing, 5034, 5034, 0, 0, 0, 0, 1, 1),
		(drawing, 5033, 5033, 0, 0, 0, 0, 1, 1),
		(drawing, 5032, 5032, 0, 0, 0, 0, 1, 1),
		(drawing, 5031, 5031, 0, 0, 0, 0, 1, 1),
		(drawing, 5030, 5030, 0, 0, 0, 0, 1, 1),
		(drawing, 5029, 5029, 0, 0, 0, 0, 1, 1),
		(drawing, 5028, 5028, 0, 0, 0, 0, 1, 1),
		(drawing, 5027, 5027, 0, 0, 0, 0, 1, 1),
		(drawing, 5026, 5026, 0, 0, 0, 0, 1, 1),
		(drawing, 5025, 5025, 0, 0, 0, 0, 1, 1),
		(drawing, 5024, 5024, 0, 0, 0, 0, 1, 1),
		(drawing, 5023, 5023, 0, 0, 0, 0, 1, 1),
		(drawing, 5022, 5022, 0, 0, 0, 0, 1, 1),
		(drawing, 5021, 5021, 0, 0, 0, 0, 1, 1),
		(drawing, 5020, 5020, 0, 0, 0, 0, 1, 1),
		(drawing, 5019, 5019, 0, 0, 0, 0, 1, 1),
		(drawing, 5018, 5018, 0, 0, 0, 0, 1, 1),
		(drawing, 5017, 5017, 0, 0, 0, 0, 1, 1),
		(drawing, 5016, 5016, 0, 0, 0, 0, 1, 1),
		(drawing, 5015, 5015, 0, 0, 0, 0, 1, 1),
		(drawing, 5014, 5014, 0, 0, 0, 0, 1, 1),
		(drawing, 5013, 5013, 0, 0, 0, 0, 1, 1),
		(drawing, 5012, 5012, 0, 0, 0, 0, 1, 1),
		(drawing, 5011, 5011, 0, 0, 0, 0, 1, 1),
		(drawing, 5010, 5010, 0, 0, 0, 0, 1, 1),
		(drawing, 5009, 5009, 0, 0, 0, 0, 1, 1),
		(drawing, 5008, 5008, 0, 0, 0, 0, 1, 1),
		(drawing, 5007, 5007, 0, 0, 0, 0, 1, 1),
		(drawing, 5006, 5006, 0, 0, 0, 0, 1, 1),
		(drawing, 5005, 5005, 0, 0, 0, 0, 1, 1),
		(drawing, 5004, 5004, 0, 0, 0, 0, 1, 1),
		(drawing, 5003, 5003, 0, 0, 0, 0, 1, 1),
		(drawing, 5002, 5002, 0, 0, 0, 0, 1, 1),
		(drawing, 5001, 5001, 0, 0, 0, 0, 1, 1),
		(drawing, 5000, 5000, 0, 0, 0, 0, 1, 1),
		(drawing, 4999, 4999, 0, 0, 0, 0, 1, 1),
		(drawing, 4998, 4998, 0, 0, 0, 0, 1, 1),
		(drawing, 4997, 4997, 0, 0, 0, 0, 1, 1),
		(drawing, 4996, 4996, 0, 0, 0, 0, 1, 1),
		(drawing, 4995, 4995, 0, 0, 0, 0, 1, 1),
		(drawing, 4994, 4994, 0, 0, 0, 0, 1, 1),
		(drawing, 4993, 4993, 0, 0, 0, 0, 1, 1),
		(drawing, 4992, 4992, 0, 0, 0, 0, 1, 1),
		(drawing, 4991, 4991, 0, 0, 0, 0, 1, 1),
		(drawing, 4990, 4990, 0, 0, 0, 0, 1, 1),
		(drawing, 4989, 4989, 0, 0, 0, 0, 1, 1),
		(drawing, 4988, 4988, 0, 0, 0, 0, 1, 1),
		(drawing, 4987, 4987, 0, 0, 0, 0, 1, 1),
		(drawing, 4986, 4986, 0, 0, 0, 0, 1, 1),
		(drawing, 4985, 4985, 0, 0, 0, 0, 1, 1),
		(drawing, 4984, 4984, 0, 0, 0, 0, 1, 1),
		(drawing, 4983, 4983, 0, 0, 0, 0, 1, 1),
		(drawing, 4982, 4982, 0, 0, 0, 0, 1, 1),
		(drawing, 4981, 4981, 0, 0, 0, 0, 1, 1),
		(drawing, 4980, 4980, 0, 0, 0, 0, 1, 1),
		(drawing, 4979, 4979, 0, 0, 0, 0, 1, 1),
		(drawing, 4978, 4978, 0, 0, 0, 0, 1, 1),
		(drawing, 4977, 4977, 0, 0, 0, 0, 1, 1),
		(drawing, 4976, 4976, 0, 0, 0, 0, 1, 1),
		(drawing, 4975, 4975, 0, 0, 0, 0, 1, 1),
		(drawing, 4974, 4974, 0, 0, 0, 0, 1, 1),
		(drawing, 4973, 4973, 0, 0, 0, 0, 1, 1),
		(drawing, 4972, 4972, 0, 0, 0, 0, 1, 1),
		(drawing, 4971, 4971, 0, 0, 0, 0, 1, 1),
		(drawing, 4970, 4970, 0, 0, 0, 0, 1, 1),
		(drawing, 4969, 4969, 0, 0, 0, 0, 1, 1),
		(drawing, 4968, 4968, 0, 0, 0, 0, 1, 1),
		(drawing, 4967, 4967, 0, 0, 0, 0, 1, 1),
		(drawing, 4966, 4966, 0, 0, 0, 0, 1, 1),
		(drawing, 4965, 4965, 0, 0, 0, 0, 1, 1),
		(drawing, 4964, 4964, 0, 0, 0, 0, 1, 1),
		(drawing, 4963, 4963, 0, 0, 0, 0, 1, 1),
		(drawing, 4962, 4962, 0, 0, 0, 0, 1, 1),
		(drawing, 4961, 4961, 0, 0, 0, 0, 1, 1),
		(drawing, 4960, 4960, 0, 0, 0, 0, 1, 1),
		(drawing, 4959, 4959, 0, 0, 0, 0, 1, 1),
		(drawing, 4958, 4958, 0, 0, 0, 0, 1, 1),
		(drawing, 4957, 4957, 0, 0, 0, 0, 1, 1),
		(drawing, 4956, 4956, 0, 0, 0, 0, 1, 1),
		(drawing, 4955, 4955, 0, 0, 0, 0, 1, 1),
		(drawing, 4954, 4954, 0, 0, 0, 0, 1, 1),
		(drawing, 4953, 4953, 0, 0, 0, 0, 1, 1),
		(drawing, 4952, 4952, 0, 0, 0, 0, 1, 1),
		(drawing, 4951, 4951, 0, 0, 0, 0, 1, 1),
		(drawing, 4950, 4950, 0, 0, 0, 0, 1, 1),
		(drawing, 4949, 4949, 0, 0, 0, 0, 1, 1),
		(drawing, 4948, 4948, 0, 0, 0, 0, 1, 1),
		(drawing, 4947, 4947, 0, 0, 0, 0, 1, 1),
		(drawing, 4946, 4946, 0, 0, 0, 0, 1, 1),
		(drawing, 4945, 4945, 0, 0, 0, 0, 1, 1),
		(drawing, 4944, 4944, 0, 0, 0, 0, 1, 1),
		(drawing, 4943, 4943, 0, 0, 0, 0, 1, 1),
		(drawing, 4942, 4942, 0, 0, 0, 0, 1, 1),
		(drawing, 4941, 4941, 0, 0, 0, 0, 1, 1),
		(drawing, 4940, 4940, 0, 0, 0, 0, 1, 1),
		(drawing, 4939, 4939, 0, 0, 0, 0, 1, 1),
		(drawing, 4938, 4938, 0, 0, 0, 0, 1, 1),
		(drawing, 4937, 4937, 0, 0, 0, 0, 1, 1),
		(drawing, 4936, 4936, 0, 0, 0, 0, 1, 1),
		(drawing, 4935, 4935, 0, 0, 0, 0, 1, 1),
		(drawing, 4934, 4934, 0, 0, 0, 0, 1, 1),
		(drawing, 4933, 4933, 0, 0, 0, 0, 1, 1),
		(drawing, 4932, 4932, 0, 0, 0, 0, 1, 1),
		(drawing, 4931, 4931, 0, 0, 0, 0, 1, 1),
		(drawing, 4930, 4930, 0, 0, 0, 0, 1, 1),
		(drawing, 4929, 4929, 0, 0, 0, 0, 1, 1),
		(drawing, 4928, 4928, 0, 0, 0, 0, 1, 1),
		(drawing, 4927, 4927, 0, 0, 0, 0, 1, 1),
		(drawing, 4926, 4926, 0, 0, 0, 0, 1, 1),
		(drawing, 4925, 4925, 0, 0, 0, 0, 1, 1),
		(drawing, 4924, 4924, 0, 0, 0, 0, 1, 1),
		(drawing, 4923, 4923, 0, 0, 0, 0, 1, 1),
		(drawing, 4922, 4922, 0, 0, 0, 0, 1, 1),
		(drawing, 4921, 4921, 0, 0, 0, 0, 1, 1),
		(drawing, 4920, 4920, 0, 0, 0, 0, 1, 1),
		(drawing, 4919, 4919, 0, 0, 0, 0, 1, 1),
		(drawing, 4918, 4918, 0, 0, 0, 0, 1, 1),
		(drawing, 4917, 4917, 0, 0, 0, 0, 1, 1),
		(drawing, 4916, 4916, 0, 0, 0, 0, 1, 1),
		(drawing, 4915, 4915, 0, 0, 0, 0, 1, 1),
		(drawing, 4914, 4914, 0, 0, 0, 0, 1, 1),
		(drawing, 4913, 4913, 0, 0, 0, 0, 1, 1),
		(drawing, 4912, 4912, 0, 0, 0, 0, 1, 1),
		(drawing, 4911, 4911, 0, 0, 0, 0, 1, 1),
		(drawing, 4910, 4910, 0, 0, 0, 0, 1, 1),
		(drawing, 4909, 4909, 0, 0, 0, 0, 1, 1),
		(drawing, 4908, 4908, 0, 0, 0, 0, 1, 1),
		(drawing, 4907, 4907, 0, 0, 0, 0, 1, 1),
		(drawing, 4906, 4906, 0, 0, 0, 0, 1, 1),
		(drawing, 4905, 4905, 0, 0, 0, 0, 1, 1),
		(drawing, 4904, 4904, 0, 0, 0, 0, 1, 1),
		(drawing, 4903, 4903, 0, 0, 0, 0, 1, 1),
		(drawing, 4902, 4902, 0, 0, 0, 0, 1, 1),
		(drawing, 4901, 4901, 0, 0, 0, 0, 1, 1),
		(drawing, 4900, 4900, 0, 0, 0, 0, 1, 1),
		(drawing, 4899, 4899, 0, 0, 0, 0, 1, 1),
		(drawing, 4898, 4898, 0, 0, 0, 0, 1, 1),
		(drawing, 4897, 4897, 0, 0, 0, 0, 1, 1),
		(drawing, 4896, 4896, 0, 0, 0, 0, 1, 1),
		(drawing, 4895, 4895, 0, 0, 0, 0, 1, 1),
		(drawing, 4894, 4894, 0, 0, 0, 0, 1, 1),
		(drawing, 4893, 4893, 0, 0, 0, 0, 1, 1),
		(drawing, 4892, 4892, 0, 0, 0, 0, 1, 1),
		(drawing, 4891, 4891, 0, 0, 0, 0, 1, 1),
		(drawing, 4890, 4890, 0, 0, 0, 0, 1, 1),
		(drawing, 4889, 4889, 0, 0, 0, 0, 1, 1),
		(drawing, 4888, 4888, 0, 0, 0, 0, 1, 1),
		(drawing, 4887, 4887, 0, 0, 0, 0, 1, 1),
		(drawing, 4886, 4886, 0, 0, 0, 0, 1, 1),
		(drawing, 4885, 4885, 0, 0, 0, 0, 1, 1),
		(drawing, 4884, 4884, 0, 0, 0, 0, 1, 1),
		(drawing, 4883, 4883, 0, 0, 0, 0, 1, 1),
		(drawing, 4882, 4882, 0, 0, 0, 0, 1, 1),
		(drawing, 4881, 4881, 0, 0, 0, 0, 1, 1),
		(drawing, 4880, 4880, 0, 0, 0, 0, 1, 1),
		(drawing, 4879, 4879, 0, 0, 0, 0, 1, 1),
		(drawing, 4878, 4878, 0, 0, 0, 0, 1, 1),
		(drawing, 4877, 4877, 0, 0, 0, 0, 1, 1),
		(drawing, 4876, 4876, 0, 0, 0, 0, 1, 1),
		(drawing, 4875, 4875, 0, 0, 0, 0, 1, 1),
		(drawing, 4874, 4874, 0, 0, 0, 0, 1, 1),
		(drawing, 4873, 4873, 0, 0, 0, 0, 1, 1),
		(drawing, 4872, 4872, 0, 0, 0, 0, 1, 1),
		(drawing, 4871, 4871, 0, 0, 0, 0, 1, 1),
		(drawing, 4870, 4870, 0, 0, 0, 0, 1, 1),
		(drawing, 4869, 4869, 0, 0, 0, 0, 1, 1),
		(drawing, 4868, 4868, 0, 0, 0, 0, 1, 1),
		(drawing, 4867, 4867, 0, 0, 0, 0, 1, 1),
		(drawing, 4866, 4866, 0, 0, 0, 0, 1, 1),
		(drawing, 4865, 4865, 0, 0, 0, 0, 1, 1),
		(drawing, 4864, 4864, 0, 0, 0, 0, 1, 1),
		(drawing, 4863, 4863, 0, 0, 0, 0, 1, 1),
		(drawing, 4862, 4862, 0, 0, 0, 0, 1, 1),
		(drawing, 4861, 4861, 0, 0, 0, 0, 1, 1),
		(drawing, 4860, 4860, 0, 0, 0, 0, 1, 1),
		(drawing, 4859, 4859, 0, 0, 0, 0, 1, 1),
		(drawing, 4858, 4858, 0, 0, 0, 0, 1, 1),
		(drawing, 4857, 4857, 0, 0, 0, 0, 1, 1),
		(drawing, 4856, 4856, 0, 0, 0, 0, 1, 1),
		(drawing, 4855, 4855, 0, 0, 0, 0, 1, 1),
		(drawing, 4854, 4854, 0, 0, 0, 0, 1, 1),
		(drawing, 4853, 4853, 0, 0, 0, 0, 1, 1),
		(drawing, 4852, 4852, 0, 0, 0, 0, 1, 1),
		(drawing, 4851, 4851, 0, 0, 0, 0, 1, 1),
		(drawing, 4850, 4850, 0, 0, 0, 0, 1, 1),
		(drawing, 4849, 4849, 0, 0, 0, 0, 1, 1),
		(drawing, 4848, 4848, 0, 0, 0, 0, 1, 1),
		(drawing, 4847, 4847, 0, 0, 0, 0, 1, 1),
		(drawing, 4846, 4846, 0, 0, 0, 0, 1, 1),
		(drawing, 4845, 4845, 0, 0, 0, 0, 1, 1),
		(drawing, 4844, 4844, 0, 0, 0, 0, 1, 1),
		(drawing, 4843, 4843, 0, 0, 0, 0, 1, 1),
		(drawing, 4842, 4842, 0, 0, 0, 0, 1, 1),
		(drawing, 4841, 4841, 0, 0, 0, 0, 1, 1),
		(drawing, 4840, 4840, 0, 0, 0, 0, 1, 1),
		(drawing, 4839, 4839, 0, 0, 0, 0, 1, 1),
		(drawing, 4838, 4838, 0, 0, 0, 0, 1, 1),
		(drawing, 4837, 4837, 0, 0, 0, 0, 1, 1),
		(drawing, 4836, 4836, 0, 0, 0, 0, 1, 1),
		(drawing, 4835, 4835, 0, 0, 0, 0, 1, 1),
		(drawing, 4834, 4834, 0, 0, 0, 0, 1, 1),
		(drawing, 4833, 4833, 0, 0, 0, 0, 1, 1),
		(drawing, 4832, 4832, 0, 0, 0, 0, 1, 1),
		(drawing, 4831, 4831, 0, 0, 0, 0, 1, 1),
		(drawing, 4830, 4830, 0, 0, 0, 0, 1, 1),
		(drawing, 4829, 4829, 0, 0, 0, 0, 1, 1),
		(drawing, 4828, 4828, 0, 0, 0, 0, 1, 1),
		(drawing, 4827, 4827, 0, 0, 0, 0, 1, 1),
		(drawing, 4826, 4826, 0, 0, 0, 0, 1, 1),
		(drawing, 4825, 4825, 0, 0, 0, 0, 1, 1),
		(drawing, 4824, 4824, 0, 0, 0, 0, 1, 1),
		(drawing, 4823, 4823, 0, 0, 0, 0, 1, 1),
		(drawing, 4822, 4822, 0, 0, 0, 0, 1, 1),
		(drawing, 4821, 4821, 0, 0, 0, 0, 1, 1),
		(drawing, 4820, 4820, 0, 0, 0, 0, 1, 1),
		(drawing, 4819, 4819, 0, 0, 0, 0, 1, 1),
		(drawing, 4818, 4818, 0, 0, 0, 0, 1, 1),
		(drawing, 4817, 4817, 0, 0, 0, 0, 1, 1),
		(drawing, 4816, 4816, 0, 0, 0, 0, 1, 1),
		(drawing, 4815, 4815, 0, 0, 0, 0, 1, 1),
		(drawing, 4814, 4814, 0, 0, 0, 0, 1, 1),
		(drawing, 4813, 4813, 0, 0, 0, 0, 1, 1),
		(drawing, 4812, 4812, 0, 0, 0, 0, 1, 1),
		(drawing, 4811, 4811, 0, 0, 0, 0, 1, 1),
		(drawing, 4810, 4810, 0, 0, 0, 0, 1, 1),
		(drawing, 4809, 4809, 0, 0, 0, 0, 1, 1),
		(drawing, 4808, 4808, 0, 0, 0, 0, 1, 1),
		(drawing, 4807, 4807, 0, 0, 0, 0, 1, 1),
		(drawing, 4806, 4806, 0, 0, 0, 0, 1, 1),
		(drawing, 4805, 4805, 0, 0, 0, 0, 1, 1),
		(drawing, 4804, 4804, 0, 0, 0, 0, 1, 1),
		(drawing, 4803, 4803, 0, 0, 0, 0, 1, 1),
		(drawing, 4802, 4802, 0, 0, 0, 0, 1, 1),
		(drawing, 4801, 4801, 0, 0, 0, 0, 1, 1),
		(drawing, 4800, 4800, 0, 0, 0, 0, 1, 1),
		(drawing, 4799, 4799, 0, 0, 0, 0, 1, 1),
		(drawing, 4798, 4798, 0, 0, 0, 0, 1, 1),
		(drawing, 4797, 4797, 0, 0, 0, 0, 1, 1),
		(drawing, 4796, 4796, 0, 0, 0, 0, 1, 1),
		(drawing, 4795, 4795, 0, 0, 0, 0, 1, 1),
		(drawing, 4794, 4794, 0, 0, 0, 0, 1, 1),
		(drawing, 4793, 4793, 0, 0, 0, 0, 1, 1),
		(drawing, 4792, 4792, 0, 0, 0, 0, 1, 1),
		(drawing, 4791, 4791, 0, 0, 0, 0, 1, 1),
		(drawing, 4790, 4790, 0, 0, 0, 0, 1, 1),
		(drawing, 4789, 4789, 0, 0, 0, 0, 1, 1),
		(drawing, 4788, 4788, 0, 0, 0, 0, 1, 1),
		(drawing, 4787, 4787, 0, 0, 0, 0, 1, 1),
		(drawing, 4786, 4786, 0, 0, 0, 0, 1, 1),
		(drawing, 4785, 4785, 0, 0, 0, 0, 1, 1),
		(drawing, 4784, 4784, 0, 0, 0, 0, 1, 1),
		(drawing, 4783, 4783, 0, 0, 0, 0, 1, 1),
		(drawing, 4782, 4782, 0, 0, 0, 0, 1, 1),
		(drawing, 4781, 4781, 0, 0, 0, 0, 1, 1),
		(drawing, 4780, 4780, 0, 0, 0, 0, 1, 1),
		(drawing, 4779, 4779, 0, 0, 0, 0, 1, 1),
		(drawing, 4778, 4778, 0, 0, 0, 0, 1, 1),
		(drawing, 4777, 4777, 0, 0, 0, 0, 1, 1),
		(drawing, 4776, 4776, 0, 0, 0, 0, 1, 1),
		(drawing, 4775, 4775, 0, 0, 0, 0, 1, 1),
		(drawing, 4774, 4774, 0, 0, 0, 0, 1, 1),
		(drawing, 4773, 4773, 0, 0, 0, 0, 1, 1),
		(drawing, 4772, 4772, 0, 0, 0, 0, 1, 1),
		(drawing, 4771, 4771, 0, 0, 0, 0, 1, 1),
		(drawing, 4770, 4770, 0, 0, 0, 0, 1, 1),
		(drawing, 4769, 4769, 0, 0, 0, 0, 1, 1),
		(drawing, 4768, 4768, 0, 0, 0, 0, 1, 1),
		(drawing, 4767, 4767, 0, 0, 0, 0, 1, 1),
		(drawing, 4766, 4766, 0, 0, 0, 0, 1, 1),
		(drawing, 4765, 4765, 0, 0, 0, 0, 1, 1),
		(drawing, 4764, 4764, 0, 0, 0, 0, 1, 1),
		(drawing, 4763, 4763, 0, 0, 0, 0, 1, 1),
		(drawing, 4762, 4762, 0, 0, 0, 0, 1, 1),
		(drawing, 4761, 4761, 0, 0, 0, 0, 1, 1),
		(drawing, 4760, 4760, 0, 0, 0, 0, 1, 1),
		(drawing, 4759, 4759, 0, 0, 0, 0, 1, 1),
		(drawing, 4758, 4758, 0, 0, 0, 0, 1, 1),
		(drawing, 4757, 4757, 0, 0, 0, 0, 1, 1),
		(drawing, 4756, 4756, 0, 0, 0, 0, 1, 1),
		(drawing, 4755, 4755, 0, 0, 0, 0, 1, 1),
		(drawing, 4754, 4754, 0, 0, 0, 0, 1, 1),
		(drawing, 4753, 4753, 0, 0, 0, 0, 1, 1),
		(drawing, 4752, 4752, 0, 0, 0, 0, 1, 1),
		(drawing, 4751, 4751, 0, 0, 0, 0, 1, 1),
		(drawing, 4750, 4750, 0, 0, 0, 0, 1, 1),
		(drawing, 4749, 4749, 0, 0, 0, 0, 1, 1),
		(drawing, 4748, 4748, 0, 0, 0, 0, 1, 1),
		(drawing, 4747, 4747, 0, 0, 0, 0, 1, 1),
		(drawing, 4746, 4746, 0, 0, 0, 0, 1, 1),
		(drawing, 4745, 4745, 0, 0, 0, 0, 1, 1),
		(drawing, 4744, 4744, 0, 0, 0, 0, 1, 1),
		(drawing, 4743, 4743, 0, 0, 0, 0, 1, 1),
		(drawing, 4742, 4742, 0, 0, 0, 0, 1, 1),
		(drawing, 4741, 4741, 0, 0, 0, 0, 1, 1),
		(drawing, 4740, 4740, 0, 0, 0, 0, 1, 1),
		(drawing, 4739, 4739, 0, 0, 0, 0, 1, 1),
		(drawing, 4738, 4738, 0, 0, 0, 0, 1, 1),
		(drawing, 4737, 4737, 0, 0, 0, 0, 1, 1),
		(drawing, 4736, 4736, 0, 0, 0, 0, 1, 1),
		(drawing, 4735, 4735, 0, 0, 0, 0, 1, 1),
		(drawing, 4734, 4734, 0, 0, 0, 0, 1, 1),
		(drawing, 4733, 4733, 0, 0, 0, 0, 1, 1),
		(drawing, 4732, 4732, 0, 0, 0, 0, 1, 1),
		(drawing, 4731, 4731, 0, 0, 0, 0, 1, 1),
		(drawing, 4730, 4730, 0, 0, 0, 0, 1, 1),
		(drawing, 4729, 4729, 0, 0, 0, 0, 1, 1),
		(drawing, 4728, 4728, 0, 0, 0, 0, 1, 1),
		(drawing, 4727, 4727, 0, 0, 0, 0, 1, 1),
		(drawing, 4726, 4726, 0, 0, 0, 0, 1, 1),
		(drawing, 4725, 4725, 0, 0, 0, 0, 1, 1),
		(drawing, 4724, 4724, 0, 0, 0, 0, 1, 1),
		(drawing, 4723, 4723, 0, 0, 0, 0, 1, 1),
		(drawing, 4722, 4722, 0, 0, 0, 0, 1, 1),
		(drawing, 4721, 4721, 0, 0, 0, 0, 1, 1),
		(drawing, 4720, 4720, 0, 0, 0, 0, 1, 1),
		(drawing, 4719, 4719, 0, 0, 0, 0, 1, 1),
		(drawing, 4718, 4718, 0, 0, 0, 0, 1, 1),
		(drawing, 4717, 4717, 0, 0, 0, 0, 1, 1),
		(drawing, 4716, 4716, 0, 0, 0, 0, 1, 1),
		(drawing, 4715, 4715, 0, 0, 0, 0, 1, 1),
		(drawing, 4714, 4714, 0, 0, 0, 0, 1, 1),
		(drawing, 4713, 4713, 0, 0, 0, 0, 1, 1),
		(drawing, 4712, 4712, 0, 0, 0, 0, 1, 1),
		(drawing, 4711, 4711, 0, 0, 0, 0, 1, 1),
		(drawing, 4710, 4710, 0, 0, 0, 0, 1, 1),
		(drawing, 4709, 4709, 0, 0, 0, 0, 1, 1),
		(drawing, 4708, 4708, 0, 0, 0, 0, 1, 1),
		(drawing, 4707, 4707, 0, 0, 0, 0, 1, 1),
		(drawing, 4706, 4706, 0, 0, 0, 0, 1, 1),
		(drawing, 4705, 4705, 0, 0, 0, 0, 1, 1),
		(drawing, 4704, 4704, 0, 0, 0, 0, 1, 1),
		(drawing, 4703, 4703, 0, 0, 0, 0, 1, 1),
		(drawing, 4702, 4702, 0, 0, 0, 0, 1, 1),
		(drawing, 4701, 4701, 0, 0, 0, 0, 1, 1),
		(drawing, 4700, 4700, 0, 0, 0, 0, 1, 1),
		(drawing, 4699, 4699, 0, 0, 0, 0, 1, 1),
		(drawing, 4698, 4698, 0, 0, 0, 0, 1, 1),
		(drawing, 4697, 4697, 0, 0, 0, 0, 1, 1),
		(drawing, 4696, 4696, 0, 0, 0, 0, 1, 1),
		(drawing, 4695, 4695, 0, 0, 0, 0, 1, 1),
		(drawing, 4694, 4694, 0, 0, 0, 0, 1, 1),
		(drawing, 4693, 4693, 0, 0, 0, 0, 1, 1),
		(drawing, 4692, 4692, 0, 0, 0, 0, 1, 1),
		(drawing, 4691, 4691, 0, 0, 0, 0, 1, 1),
		(drawing, 4690, 4690, 0, 0, 0, 0, 1, 1),
		(drawing, 4689, 4689, 0, 0, 0, 0, 1, 1),
		(drawing, 4688, 4688, 0, 0, 0, 0, 1, 1),
		(drawing, 4687, 4687, 0, 0, 0, 0, 1, 1),
		(drawing, 4686, 4686, 0, 0, 0, 0, 1, 1),
		(drawing, 4685, 4685, 0, 0, 0, 0, 1, 1),
		(drawing, 4684, 4684, 0, 0, 0, 0, 1, 1),
		(drawing, 4683, 4683, 0, 0, 0, 0, 1, 1),
		(drawing, 4682, 4682, 0, 0, 0, 0, 1, 1),
		(drawing, 4681, 4681, 0, 0, 0, 0, 1, 1),
		(drawing, 4680, 4680, 0, 0, 0, 0, 1, 1),
		(drawing, 4679, 4679, 0, 0, 0, 0, 1, 1),
		(drawing, 4678, 4678, 0, 0, 0, 0, 1, 1),
		(drawing, 4677, 4677, 0, 0, 0, 0, 1, 1),
		(drawing, 4676, 4676, 0, 0, 0, 0, 1, 1),
		(drawing, 4675, 4675, 0, 0, 0, 0, 1, 1),
		(drawing, 4674, 4674, 0, 0, 0, 0, 1, 1),
		(drawing, 4673, 4673, 0, 0, 0, 0, 1, 1),
		(drawing, 4672, 4672, 0, 0, 0, 0, 1, 1),
		(drawing, 4671, 4671, 0, 0, 0, 0, 1, 1),
		(drawing, 4670, 4670, 0, 0, 0, 0, 1, 1),
		(drawing, 4669, 4669, 0, 0, 0, 0, 1, 1),
		(drawing, 4668, 4668, 0, 0, 0, 0, 1, 1),
		(drawing, 4667, 4667, 0, 0, 0, 0, 1, 1),
		(drawing, 4666, 4666, 0, 0, 0, 0, 1, 1),
		(drawing, 4665, 4665, 0, 0, 0, 0, 1, 1),
		(drawing, 4664, 4664, 0, 0, 0, 0, 1, 1),
		(drawing, 4663, 4663, 0, 0, 0, 0, 1, 1),
		(drawing, 4662, 4662, 0, 0, 0, 0, 1, 1),
		(drawing, 4661, 4661, 0, 0, 0, 0, 1, 1),
		(drawing, 4660, 4660, 0, 0, 0, 0, 1, 1),
		(drawing, 4659, 4659, 0, 0, 0, 0, 1, 1),
		(drawing, 4658, 4658, 0, 0, 0, 0, 1, 1),
		(drawing, 4657, 4657, 0, 0, 0, 0, 1, 1),
		(drawing, 4656, 4656, 0, 0, 0, 0, 1, 1),
		(drawing, 4655, 4655, 0, 0, 0, 0, 1, 1),
		(drawing, 4654, 4654, 0, 0, 0, 0, 1, 1),
		(drawing, 4653, 4653, 0, 0, 0, 0, 1, 1),
		(drawing, 4652, 4652, 0, 0, 0, 0, 1, 1),
		(drawing, 4651, 4651, 0, 0, 0, 0, 1, 1),
		(drawing, 4650, 4650, 0, 0, 0, 0, 1, 1),
		(drawing, 4649, 4649, 0, 0, 0, 0, 1, 1),
		(drawing, 4648, 4648, 0, 0, 0, 0, 1, 1),
		(drawing, 4647, 4647, 0, 0, 0, 0, 1, 1),
		(drawing, 4646, 4646, 0, 0, 0, 0, 1, 1),
		(drawing, 4645, 4645, 0, 0, 0, 0, 1, 1),
		(drawing, 4644, 4644, 0, 0, 0, 0, 1, 1),
		(drawing, 4643, 4643, 0, 0, 0, 0, 1, 1),
		(drawing, 4642, 4642, 0, 0, 0, 0, 1, 1),
		(drawing, 4641, 4641, 0, 0, 0, 0, 1, 1),
		(drawing, 4640, 4640, 0, 0, 0, 0, 1, 1),
		(drawing, 4639, 4639, 0, 0, 0, 0, 1, 1),
		(drawing, 4638, 4638, 0, 0, 0, 0, 1, 1),
		(drawing, 4637, 4637, 0, 0, 0, 0, 1, 1),
		(drawing, 4636, 4636, 0, 0, 0, 0, 1, 1),
		(drawing, 4635, 4635, 0, 0, 0, 0, 1, 1),
		(drawing, 4634, 4634, 0, 0, 0, 0, 1, 1),
		(drawing, 4633, 4633, 0, 0, 0, 0, 1, 1),
		(drawing, 4632, 4632, 0, 0, 0, 0, 1, 1),
		(drawing, 4631, 4631, 0, 0, 0, 0, 1, 1),
		(drawing, 4630, 4630, 0, 0, 0, 0, 1, 1),
		(drawing, 4629, 4629, 0, 0, 0, 0, 1, 1),
		(drawing, 4628, 4628, 0, 0, 0, 0, 1, 1),
		(drawing, 4627, 4627, 0, 0, 0, 0, 1, 1),
		(drawing, 4626, 4626, 0, 0, 0, 0, 1, 1),
		(drawing, 4625, 4625, 0, 0, 0, 0, 1, 1),
		(drawing, 4624, 4624, 0, 0, 0, 0, 1, 1),
		(drawing, 4623, 4623, 0, 0, 0, 0, 1, 1),
		(drawing, 4622, 4622, 0, 0, 0, 0, 1, 1),
		(drawing, 4621, 4621, 0, 0, 0, 0, 1, 1),
		(drawing, 4620, 4620, 0, 0, 0, 0, 1, 1),
		(drawing, 4619, 4619, 0, 0, 0, 0, 1, 1),
		(drawing, 4618, 4618, 0, 0, 0, 0, 1, 1),
		(drawing, 4617, 4617, 0, 0, 0, 0, 1, 1),
		(drawing, 4616, 4616, 0, 0, 0, 0, 1, 1),
		(drawing, 4615, 4615, 0, 0, 0, 0, 1, 1),
		(drawing, 4614, 4614, 0, 0, 0, 0, 1, 1),
		(drawing, 4613, 4613, 0, 0, 0, 0, 1, 1),
		(drawing, 4612, 4612, 0, 0, 0, 0, 1, 1),
		(drawing, 4611, 4611, 0, 0, 0, 0, 1, 1),
		(drawing, 4610, 4610, 0, 0, 0, 0, 1, 1),
		(drawing, 4609, 4609, 0, 0, 0, 0, 1, 1),
		(drawing, 4608, 4608, 0, 0, 0, 0, 1, 1),
		(drawing, 4607, 4607, 0, 0, 0, 0, 1, 1),
		(drawing, 4606, 4606, 0, 0, 0, 0, 1, 1),
		(drawing, 4605, 4605, 0, 0, 0, 0, 1, 1),
		(drawing, 4604, 4604, 0, 0, 0, 0, 1, 1),
		(drawing, 4603, 4603, 0, 0, 0, 0, 1, 1),
		(drawing, 4602, 4602, 0, 0, 0, 0, 1, 1),
		(drawing, 4601, 4601, 0, 0, 0, 0, 1, 1),
		(drawing, 4600, 4600, 0, 0, 0, 0, 1, 1),
		(drawing, 4599, 4599, 0, 0, 0, 0, 1, 1),
		(drawing, 4598, 4598, 0, 0, 0, 0, 1, 1),
		(drawing, 4597, 4597, 0, 0, 0, 0, 1, 1),
		(drawing, 4596, 4596, 0, 0, 0, 0, 1, 1),
		(drawing, 4595, 4595, 0, 0, 0, 0, 1, 1),
		(drawing, 4594, 4594, 0, 0, 0, 0, 1, 1),
		(drawing, 4593, 4593, 0, 0, 0, 0, 1, 1),
		(drawing, 4592, 4592, 0, 0, 0, 0, 1, 1),
		(drawing, 4591, 4591, 0, 0, 0, 0, 1, 1),
		(drawing, 4590, 4590, 0, 0, 0, 0, 1, 1),
		(drawing, 4589, 4589, 0, 0, 0, 0, 1, 1),
		(drawing, 4588, 4588, 0, 0, 0, 0, 1, 1),
		(drawing, 4587, 4587, 0, 0, 0, 0, 1, 1),
		(drawing, 4586, 4586, 0, 0, 0, 0, 1, 1),
		(drawing, 4585, 4585, 0, 0, 0, 0, 1, 1),
		(drawing, 4584, 4584, 0, 0, 0, 0, 1, 1),
		(drawing, 4583, 4583, 0, 0, 0, 0, 1, 1),
		(drawing, 4582, 4582, 0, 0, 0, 0, 1, 1),
		(drawing, 4581, 4581, 0, 0, 0, 0, 1, 1),
		(drawing, 4580, 4580, 0, 0, 0, 0, 1, 1),
		(drawing, 4579, 4579, 0, 0, 0, 0, 1, 1),
		(drawing, 4578, 4578, 0, 0, 0, 0, 1, 1),
		(drawing, 4577, 4577, 0, 0, 0, 0, 1, 1),
		(drawing, 4576, 4576, 0, 0, 0, 0, 1, 1),
		(drawing, 4575, 4575, 0, 0, 0, 0, 1, 1),
		(drawing, 4574, 4574, 0, 0, 0, 0, 1, 1),
		(drawing, 4573, 4573, 0, 0, 0, 0, 1, 1),
		(drawing, 4572, 4572, 0, 0, 0, 0, 1, 1),
		(drawing, 4571, 4571, 0, 0, 0, 0, 1, 1),
		(drawing, 4570, 4570, 0, 0, 0, 0, 1, 1),
		(drawing, 4569, 4569, 0, 0, 0, 0, 1, 1),
		(drawing, 4568, 4568, 0, 0, 0, 0, 1, 1),
		(drawing, 4567, 4567, 0, 0, 0, 0, 1, 1),
		(drawing, 4566, 4566, 0, 0, 0, 0, 1, 1),
		(drawing, 4565, 4565, 0, 0, 0, 0, 1, 1),
		(drawing, 4564, 4564, 0, 0, 0, 0, 1, 1),
		(drawing, 4563, 4563, 0, 0, 0, 0, 1, 1),
		(drawing, 4562, 4562, 0, 0, 0, 0, 1, 1),
		(drawing, 4561, 4561, 0, 0, 0, 0, 1, 1),
		(drawing, 4560, 4560, 0, 0, 0, 0, 1, 1),
		(drawing, 4559, 4559, 0, 0, 0, 0, 1, 1),
		(drawing, 4558, 4558, 0, 0, 0, 0, 1, 1),
		(drawing, 4557, 4557, 0, 0, 0, 0, 1, 1),
		(drawing, 4556, 4556, 0, 0, 0, 0, 1, 1),
		(drawing, 4555, 4555, 0, 0, 0, 0, 1, 1),
		(drawing, 4554, 4554, 0, 0, 0, 0, 1, 1),
		(drawing, 4553, 4553, 0, 0, 0, 0, 1, 1),
		(drawing, 4552, 4552, 0, 0, 0, 0, 1, 1),
		(drawing, 4551, 4551, 0, 0, 0, 0, 1, 1),
		(drawing, 4550, 4550, 0, 0, 0, 0, 1, 1),
		(drawing, 4549, 4549, 0, 0, 0, 0, 1, 1),
		(drawing, 4548, 4548, 0, 0, 0, 0, 1, 1),
		(drawing, 4547, 4547, 0, 0, 0, 0, 1, 1),
		(drawing, 4546, 4546, 0, 0, 0, 0, 1, 1),
		(drawing, 4545, 4545, 0, 0, 0, 0, 1, 1),
		(drawing, 4544, 4544, 0, 0, 0, 0, 1, 1),
		(drawing, 4543, 4543, 0, 0, 0, 0, 1, 1),
		(drawing, 4542, 4542, 0, 0, 0, 0, 1, 1),
		(drawing, 4541, 4541, 0, 0, 0, 0, 1, 1),
		(drawing, 4540, 4540, 0, 0, 0, 0, 1, 1),
		(drawing, 4539, 4539, 0, 0, 0, 0, 1, 1),
		(drawing, 4538, 4538, 0, 0, 0, 0, 1, 1),
		(drawing, 4537, 4537, 0, 0, 0, 0, 1, 1),
		(drawing, 4536, 4536, 0, 0, 0, 0, 1, 1),
		(drawing, 4535, 4535, 0, 0, 0, 0, 1, 1),
		(drawing, 4534, 4534, 0, 0, 0, 0, 1, 1),
		(drawing, 4533, 4533, 0, 0, 0, 0, 1, 1),
		(drawing, 4532, 4532, 0, 0, 0, 0, 1, 1),
		(drawing, 4531, 4531, 0, 0, 0, 0, 1, 1),
		(drawing, 4530, 4530, 0, 0, 0, 0, 1, 1),
		(drawing, 4529, 4529, 0, 0, 0, 0, 1, 1),
		(drawing, 4528, 4528, 0, 0, 0, 0, 1, 1),
		(drawing, 4527, 4527, 0, 0, 0, 0, 1, 1),
		(drawing, 4526, 4526, 0, 0, 0, 0, 1, 1),
		(drawing, 4525, 4525, 0, 0, 0, 0, 1, 1),
		(drawing, 4524, 4524, 0, 0, 0, 0, 1, 1),
		(drawing, 4523, 4523, 0, 0, 0, 0, 1, 1),
		(drawing, 4522, 4522, 0, 0, 0, 0, 1, 1),
		(drawing, 4521, 4521, 0, 0, 0, 0, 1, 1),
		(drawing, 4520, 4520, 0, 0, 0, 0, 1, 1),
		(drawing, 4519, 4519, 0, 0, 0, 0, 1, 1),
		(drawing, 4518, 4518, 0, 0, 0, 0, 1, 1),
		(drawing, 4517, 4517, 0, 0, 0, 0, 1, 1),
		(drawing, 4516, 4516, 0, 0, 0, 0, 1, 1),
		(drawing, 4515, 4515, 0, 0, 0, 0, 1, 1),
		(drawing, 4514, 4514, 0, 0, 0, 0, 1, 1),
		(drawing, 4513, 4513, 0, 0, 0, 0, 1, 1),
		(drawing, 4512, 4512, 0, 0, 0, 0, 1, 1),
		(drawing, 4511, 4511, 0, 0, 0, 0, 1, 1),
		(drawing, 4510, 4510, 0, 0, 0, 0, 1, 1),
		(drawing, 4509, 4509, 0, 0, 0, 0, 1, 1),
		(drawing, 4508, 4508, 0, 0, 0, 0, 1, 1),
		(drawing, 4507, 4507, 0, 0, 0, 0, 1, 1),
		(drawing, 4506, 4506, 0, 0, 0, 0, 1, 1),
		(drawing, 4505, 4505, 0, 0, 0, 0, 1, 1),
		(drawing, 4504, 4504, 0, 0, 0, 0, 1, 1),
		(drawing, 4503, 4503, 0, 0, 0, 0, 1, 1),
		(drawing, 4502, 4502, 0, 0, 0, 0, 1, 1),
		(drawing, 4501, 4501, 0, 0, 0, 0, 1, 1),
		(drawing, 4500, 4500, 0, 0, 0, 0, 1, 1),
		(drawing, 4499, 4499, 0, 0, 0, 0, 1, 1),
		(drawing, 4498, 4498, 0, 0, 0, 0, 1, 1),
		(drawing, 4497, 4497, 0, 0, 0, 0, 1, 1),
		(drawing, 4496, 4496, 0, 0, 0, 0, 1, 1),
		(drawing, 4495, 4495, 0, 0, 0, 0, 1, 1),
		(drawing, 4494, 4494, 0, 0, 0, 0, 1, 1),
		(drawing, 4493, 4493, 0, 0, 0, 0, 1, 1),
		(drawing, 4492, 4492, 0, 0, 0, 0, 1, 1),
		(drawing, 4491, 4491, 0, 0, 0, 0, 1, 1),
		(drawing, 4490, 4490, 0, 0, 0, 0, 1, 1),
		(drawing, 4489, 4489, 0, 0, 0, 0, 1, 1),
		(drawing, 4488, 4488, 0, 0, 0, 0, 1, 1),
		(drawing, 4487, 4487, 0, 0, 0, 0, 1, 1),
		(drawing, 4486, 4486, 0, 0, 0, 0, 1, 1),
		(drawing, 4485, 4485, 0, 0, 0, 0, 1, 1),
		(drawing, 4484, 4484, 0, 0, 0, 0, 1, 1),
		(drawing, 4483, 4483, 0, 0, 0, 0, 1, 1),
		(drawing, 4482, 4482, 0, 0, 0, 0, 1, 1),
		(drawing, 4481, 4481, 0, 0, 0, 0, 1, 1),
		(drawing, 4480, 4480, 0, 0, 0, 0, 1, 1),
		(drawing, 4479, 4479, 0, 0, 0, 0, 1, 1),
		(drawing, 4478, 4478, 0, 0, 0, 0, 1, 1),
		(drawing, 4477, 4477, 0, 0, 0, 0, 1, 1),
		(drawing, 4476, 4476, 0, 0, 0, 0, 1, 1),
		(drawing, 4475, 4475, 0, 0, 0, 0, 1, 1),
		(drawing, 4474, 4474, 0, 0, 0, 0, 1, 1),
		(drawing, 4473, 4473, 0, 0, 0, 0, 1, 1),
		(drawing, 4472, 4472, 0, 0, 0, 0, 1, 1),
		(drawing, 4471, 4471, 0, 0, 0, 0, 1, 1),
		(drawing, 4470, 4470, 0, 0, 0, 0, 1, 1),
		(drawing, 4469, 4469, 0, 0, 0, 0, 1, 1),
		(drawing, 4468, 4468, 0, 0, 0, 0, 1, 1),
		(drawing, 4467, 4467, 0, 0, 0, 0, 1, 1),
		(drawing, 4466, 4466, 0, 0, 0, 0, 1, 1),
		(drawing, 4465, 4465, 0, 0, 0, 0, 1, 1),
		(drawing, 4464, 4464, 0, 0, 0, 0, 1, 1),
		(drawing, 4463, 4463, 0, 0, 0, 0, 1, 1),
		(drawing, 4462, 4462, 0, 0, 0, 0, 1, 1),
		(drawing, 4461, 4461, 0, 0, 0, 0, 1, 1),
		(drawing, 4460, 4460, 0, 0, 0, 0, 1, 1),
		(drawing, 4459, 4459, 0, 0, 0, 0, 1, 1),
		(drawing, 4458, 4458, 0, 0, 0, 0, 1, 1),
		(drawing, 4457, 4457, 0, 0, 0, 0, 1, 1),
		(drawing, 4456, 4456, 0, 0, 0, 0, 1, 1),
		(drawing, 4455, 4455, 0, 0, 0, 0, 1, 1),
		(drawing, 4454, 4454, 0, 0, 0, 0, 1, 1),
		(drawing, 4453, 4453, 0, 0, 0, 0, 1, 1),
		(drawing, 4452, 4452, 0, 0, 0, 0, 1, 1),
		(drawing, 4451, 4451, 0, 0, 0, 0, 1, 1),
		(drawing, 4450, 4450, 0, 0, 0, 0, 1, 1),
		(drawing, 4449, 4449, 0, 0, 0, 0, 1, 1),
		(drawing, 4448, 4448, 0, 0, 0, 0, 1, 1),
		(drawing, 4447, 4447, 0, 0, 0, 0, 1, 1),
		(drawing, 4446, 4446, 0, 0, 0, 0, 1, 1),
		(drawing, 4445, 4445, 0, 0, 0, 0, 1, 1),
		(drawing, 4444, 4444, 0, 0, 0, 0, 1, 1),
		(drawing, 4443, 4443, 0, 0, 0, 0, 1, 1),
		(drawing, 4442, 4442, 0, 0, 0, 0, 1, 1),
		(drawing, 4441, 4441, 0, 0, 0, 0, 1, 1),
		(drawing, 4440, 4440, 0, 0, 0, 0, 1, 1),
		(drawing, 4439, 4439, 0, 0, 0, 0, 1, 1),
		(drawing, 4438, 4438, 0, 0, 0, 0, 1, 1),
		(drawing, 4437, 4437, 0, 0, 0, 0, 1, 1),
		(drawing, 4436, 4436, 0, 0, 0, 0, 1, 1),
		(drawing, 4435, 4435, 0, 0, 0, 0, 1, 1),
		(drawing, 4434, 4434, 0, 0, 0, 0, 1, 1),
		(drawing, 4433, 4433, 0, 0, 0, 0, 1, 1),
		(drawing, 4432, 4432, 0, 0, 0, 0, 1, 1),
		(drawing, 4431, 4431, 0, 0, 0, 0, 1, 1),
		(drawing, 4430, 4430, 0, 0, 0, 0, 1, 1),
		(drawing, 4429, 4429, 0, 0, 0, 0, 1, 1),
		(drawing, 4428, 4428, 0, 0, 0, 0, 1, 1),
		(drawing, 4427, 4427, 0, 0, 0, 0, 1, 1),
		(drawing, 4426, 4426, 0, 0, 0, 0, 1, 1),
		(drawing, 4425, 4425, 0, 0, 0, 0, 1, 1),
		(drawing, 4424, 4424, 0, 0, 0, 0, 1, 1),
		(drawing, 4423, 4423, 0, 0, 0, 0, 1, 1),
		(drawing, 4422, 4422, 0, 0, 0, 0, 1, 1),
		(drawing, 4421, 4421, 0, 0, 0, 0, 1, 1),
		(drawing, 4420, 4420, 0, 0, 0, 0, 1, 1),
		(drawing, 4419, 4419, 0, 0, 0, 0, 1, 1),
		(drawing, 4418, 4418, 0, 0, 0, 0, 1, 1),
		(drawing, 4417, 4417, 0, 0, 0, 0, 1, 1),
		(drawing, 4416, 4416, 0, 0, 0, 0, 1, 1),
		(drawing, 4415, 4415, 0, 0, 0, 0, 1, 1),
		(drawing, 4414, 4414, 0, 0, 0, 0, 1, 1),
		(drawing, 4413, 4413, 0, 0, 0, 0, 1, 1),
		(drawing, 4412, 4412, 0, 0, 0, 0, 1, 1),
		(drawing, 4411, 4411, 0, 0, 0, 0, 1, 1),
		(drawing, 4410, 4410, 0, 0, 0, 0, 1, 1),
		(drawing, 4409, 4409, 0, 0, 0, 0, 1, 1),
		(drawing, 4408, 4408, 0, 0, 0, 0, 1, 1),
		(drawing, 4407, 4407, 0, 0, 0, 0, 1, 1),
		(drawing, 4406, 4406, 0, 0, 0, 0, 1, 1),
		(drawing, 4405, 4405, 0, 0, 0, 0, 1, 1),
		(drawing, 4404, 4404, 0, 0, 0, 0, 1, 1),
		(drawing, 4403, 4403, 0, 0, 0, 0, 1, 1),
		(drawing, 4402, 4402, 0, 0, 0, 0, 1, 1),
		(drawing, 4401, 4401, 0, 0, 0, 0, 1, 1),
		(drawing, 4400, 4400, 0, 0, 0, 0, 1, 1),
		(drawing, 4399, 4399, 0, 0, 0, 0, 1, 1),
		(drawing, 4398, 4398, 0, 0, 0, 0, 1, 1),
		(drawing, 4397, 4397, 0, 0, 0, 0, 1, 1),
		(drawing, 4396, 4396, 0, 0, 0, 0, 1, 1),
		(drawing, 4395, 4395, 0, 0, 0, 0, 1, 1),
		(drawing, 4394, 4394, 0, 0, 0, 0, 1, 1),
		(drawing, 4393, 4393, 0, 0, 0, 0, 1, 1),
		(drawing, 4392, 4392, 0, 0, 0, 0, 1, 1),
		(drawing, 4391, 4391, 0, 0, 0, 0, 1, 1),
		(drawing, 4390, 4390, 0, 0, 0, 0, 1, 1),
		(drawing, 4389, 4389, 0, 0, 0, 0, 1, 1),
		(drawing, 4388, 4388, 0, 0, 0, 0, 1, 1),
		(drawing, 4387, 4387, 0, 0, 0, 0, 1, 1),
		(drawing, 4386, 4386, 0, 0, 0, 0, 1, 1),
		(drawing, 4385, 4385, 0, 0, 0, 0, 1, 1),
		(drawing, 4384, 4384, 0, 0, 0, 0, 1, 1),
		(drawing, 4383, 4383, 0, 0, 0, 0, 1, 1),
		(drawing, 4382, 4382, 0, 0, 0, 0, 1, 1),
		(drawing, 4381, 4381, 0, 0, 0, 0, 1, 1),
		(drawing, 4380, 4380, 0, 0, 0, 0, 1, 1),
		(drawing, 4379, 4379, 0, 0, 0, 0, 1, 1),
		(drawing, 4378, 4378, 0, 0, 0, 0, 1, 1),
		(drawing, 4377, 4377, 0, 0, 0, 0, 1, 1),
		(drawing, 4376, 4376, 0, 0, 0, 0, 1, 1),
		(drawing, 4375, 4375, 0, 0, 0, 0, 1, 1),
		(drawing, 4374, 4374, 0, 0, 0, 0, 1, 1),
		(drawing, 4373, 4373, 0, 0, 0, 0, 1, 1),
		(drawing, 4372, 4372, 0, 0, 0, 0, 1, 1),
		(drawing, 4371, 4371, 0, 0, 0, 0, 1, 1),
		(drawing, 4370, 4370, 0, 0, 0, 0, 1, 1),
		(drawing, 4369, 4369, 0, 0, 0, 0, 1, 1),
		(drawing, 4368, 4368, 0, 0, 0, 0, 1, 1),
		(drawing, 4367, 4367, 0, 0, 0, 0, 1, 1),
		(drawing, 4366, 4366, 0, 0, 0, 0, 1, 1),
		(drawing, 4365, 4365, 0, 0, 0, 0, 1, 1),
		(drawing, 4364, 4364, 0, 0, 0, 0, 1, 1),
		(drawing, 4363, 4363, 0, 0, 0, 0, 1, 1),
		(drawing, 4362, 4362, 0, 0, 0, 0, 1, 1),
		(drawing, 4361, 4361, 0, 0, 0, 0, 1, 1),
		(drawing, 4360, 4360, 0, 0, 0, 0, 1, 1),
		(drawing, 4359, 4359, 0, 0, 0, 0, 1, 1),
		(drawing, 4358, 4358, 0, 0, 0, 0, 1, 1),
		(drawing, 4357, 4357, 0, 0, 0, 0, 1, 1),
		(drawing, 4356, 4356, 0, 0, 0, 0, 1, 1),
		(drawing, 4355, 4355, 0, 0, 0, 0, 1, 1),
		(drawing, 4354, 4354, 0, 0, 0, 0, 1, 1),
		(drawing, 4353, 4353, 0, 0, 0, 0, 1, 1),
		(drawing, 4352, 4352, 0, 0, 0, 0, 1, 1),
		(drawing, 4351, 4351, 0, 0, 0, 0, 1, 1),
		(drawing, 4350, 4350, 0, 0, 0, 0, 1, 1),
		(drawing, 4349, 4349, 0, 0, 0, 0, 1, 1),
		(drawing, 4348, 4348, 0, 0, 0, 0, 1, 1),
		(drawing, 4347, 4347, 0, 0, 0, 0, 1, 1),
		(drawing, 4346, 4346, 0, 0, 0, 0, 1, 1),
		(drawing, 4345, 4345, 0, 0, 0, 0, 1, 1),
		(drawing, 4344, 4344, 0, 0, 0, 0, 1, 1),
		(drawing, 4343, 4343, 0, 0, 0, 0, 1, 1),
		(drawing, 4342, 4342, 0, 0, 0, 0, 1, 1),
		(drawing, 4341, 4341, 0, 0, 0, 0, 1, 1),
		(drawing, 4340, 4340, 0, 0, 0, 0, 1, 1),
		(drawing, 4339, 4339, 0, 0, 0, 0, 1, 1),
		(drawing, 4338, 4338, 0, 0, 0, 0, 1, 1),
		(drawing, 4337, 4337, 0, 0, 0, 0, 1, 1),
		(drawing, 4336, 4336, 0, 0, 0, 0, 1, 1),
		(drawing, 4335, 4335, 0, 0, 0, 0, 1, 1),
		(drawing, 4334, 4334, 0, 0, 0, 0, 1, 1),
		(drawing, 4333, 4333, 0, 0, 0, 0, 1, 1),
		(drawing, 4332, 4332, 0, 0, 0, 0, 1, 1),
		(drawing, 4331, 4331, 0, 0, 0, 0, 1, 1),
		(drawing, 4330, 4330, 0, 0, 0, 0, 1, 1),
		(drawing, 4329, 4329, 0, 0, 0, 0, 1, 1),
		(drawing, 4328, 4328, 0, 0, 0, 0, 1, 1),
		(drawing, 4327, 4327, 0, 0, 0, 0, 1, 1),
		(drawing, 4326, 4326, 0, 0, 0, 0, 1, 1),
		(drawing, 4325, 4325, 0, 0, 0, 0, 1, 1),
		(drawing, 4324, 4324, 0, 0, 0, 0, 1, 1),
		(drawing, 4323, 4323, 0, 0, 0, 0, 1, 1),
		(drawing, 4322, 4322, 0, 0, 0, 0, 1, 1),
		(drawing, 4321, 4321, 0, 0, 0, 0, 1, 1),
		(drawing, 4320, 4320, 0, 0, 0, 0, 1, 1),
		(drawing, 4319, 4319, 0, 0, 0, 0, 1, 1),
		(drawing, 4318, 4318, 0, 0, 0, 0, 1, 1),
		(drawing, 4317, 4317, 0, 0, 0, 0, 1, 1),
		(drawing, 4316, 4316, 0, 0, 0, 0, 1, 1),
		(drawing, 4315, 4315, 0, 0, 0, 0, 1, 1),
		(drawing, 4314, 4314, 0, 0, 0, 0, 1, 1),
		(drawing, 4313, 4313, 0, 0, 0, 0, 1, 1),
		(drawing, 4312, 4312, 0, 0, 0, 0, 1, 1),
		(drawing, 4311, 4311, 0, 0, 0, 0, 1, 1),
		(drawing, 4310, 4310, 0, 0, 0, 0, 1, 1),
		(drawing, 4309, 4309, 0, 0, 0, 0, 1, 1),
		(drawing, 4308, 4308, 0, 0, 0, 0, 1, 1),
		(drawing, 4307, 4307, 0, 0, 0, 0, 1, 1),
		(drawing, 4306, 4306, 0, 0, 0, 0, 1, 1),
		(drawing, 4305, 4305, 0, 0, 0, 0, 1, 1),
		(drawing, 4304, 4304, 0, 0, 0, 0, 1, 1),
		(drawing, 4303, 4303, 0, 0, 0, 0, 1, 1),
		(drawing, 4302, 4302, 0, 0, 0, 0, 1, 1),
		(drawing, 4301, 4301, 0, 0, 0, 0, 1, 1),
		(drawing, 4300, 4300, 0, 0, 0, 0, 1, 1),
		(drawing, 4299, 4299, 0, 0, 0, 0, 1, 1),
		(drawing, 4298, 4298, 0, 0, 0, 0, 1, 1),
		(drawing, 4297, 4297, 0, 0, 0, 0, 1, 1),
		(drawing, 4296, 4296, 0, 0, 0, 0, 1, 1),
		(drawing, 4295, 4295, 0, 0, 0, 0, 1, 1),
		(drawing, 4294, 4294, 0, 0, 0, 0, 1, 1),
		(drawing, 4293, 4293, 0, 0, 0, 0, 1, 1),
		(drawing, 4292, 4292, 0, 0, 0, 0, 1, 1),
		(drawing, 4291, 4291, 0, 0, 0, 0, 1, 1),
		(drawing, 4290, 4290, 0, 0, 0, 0, 1, 1),
		(drawing, 4289, 4289, 0, 0, 0, 0, 1, 1),
		(drawing, 4288, 4288, 0, 0, 0, 0, 1, 1),
		(drawing, 4287, 4287, 0, 0, 0, 0, 1, 1),
		(drawing, 4286, 4286, 0, 0, 0, 0, 1, 1),
		(drawing, 4285, 4285, 0, 0, 0, 0, 1, 1),
		(drawing, 4284, 4284, 0, 0, 0, 0, 1, 1),
		(drawing, 4283, 4283, 0, 0, 0, 0, 1, 1),
		(drawing, 4282, 4282, 0, 0, 0, 0, 1, 1),
		(drawing, 4281, 4281, 0, 0, 0, 0, 1, 1),
		(drawing, 4280, 4280, 0, 0, 0, 0, 1, 1),
		(drawing, 4279, 4279, 0, 0, 0, 0, 1, 1),
		(drawing, 4278, 4278, 0, 0, 0, 0, 1, 1),
		(drawing, 4277, 4277, 0, 0, 0, 0, 1, 1),
		(drawing, 4276, 4276, 0, 0, 0, 0, 1, 1),
		(drawing, 4275, 4275, 0, 0, 0, 0, 1, 1),
		(drawing, 4274, 4274, 0, 0, 0, 0, 1, 1),
		(drawing, 4273, 4273, 0, 0, 0, 0, 1, 1),
		(drawing, 4272, 4272, 0, 0, 0, 0, 1, 1),
		(drawing, 4271, 4271, 0, 0, 0, 0, 1, 1),
		(drawing, 4270, 4270, 0, 0, 0, 0, 1, 1),
		(drawing, 4269, 4269, 0, 0, 0, 0, 1, 1),
		(drawing, 4268, 4268, 0, 0, 0, 0, 1, 1),
		(drawing, 4267, 4267, 0, 0, 0, 0, 1, 1),
		(drawing, 4266, 4266, 0, 0, 0, 0, 1, 1),
		(drawing, 4265, 4265, 0, 0, 0, 0, 1, 1),
		(drawing, 4264, 4264, 0, 0, 0, 0, 1, 1),
		(drawing, 4263, 4263, 0, 0, 0, 0, 1, 1),
		(drawing, 4262, 4262, 0, 0, 0, 0, 1, 1),
		(drawing, 4261, 4261, 0, 0, 0, 0, 1, 1),
		(drawing, 4260, 4260, 0, 0, 0, 0, 1, 1),
		(drawing, 4259, 4259, 0, 0, 0, 0, 1, 1),
		(drawing, 4258, 4258, 0, 0, 0, 0, 1, 1),
		(drawing, 4257, 4257, 0, 0, 0, 0, 1, 1),
		(drawing, 4256, 4256, 0, 0, 0, 0, 1, 1),
		(drawing, 4255, 4255, 0, 0, 0, 0, 1, 1),
		(drawing, 4254, 4254, 0, 0, 0, 0, 1, 1),
		(drawing, 4253, 4253, 0, 0, 0, 0, 1, 1),
		(drawing, 4252, 4252, 0, 0, 0, 0, 1, 1),
		(drawing, 4251, 4251, 0, 0, 0, 0, 1, 1),
		(drawing, 4250, 4250, 0, 0, 0, 0, 1, 1),
		(drawing, 4249, 4249, 0, 0, 0, 0, 1, 1),
		(drawing, 4248, 4248, 0, 0, 0, 0, 1, 1),
		(drawing, 4247, 4247, 0, 0, 0, 0, 1, 1),
		(drawing, 4246, 4246, 0, 0, 0, 0, 1, 1),
		(drawing, 4245, 4245, 0, 0, 0, 0, 1, 1),
		(drawing, 4244, 4244, 0, 0, 0, 0, 1, 1),
		(drawing, 4243, 4243, 0, 0, 0, 0, 1, 1),
		(drawing, 4242, 4242, 0, 0, 0, 0, 1, 1),
		(drawing, 4241, 4241, 0, 0, 0, 0, 1, 1),
		(drawing, 4240, 4240, 0, 0, 0, 0, 1, 1),
		(drawing, 4239, 4239, 0, 0, 0, 0, 1, 1),
		(drawing, 4238, 4238, 0, 0, 0, 0, 1, 1),
		(drawing, 4237, 4237, 0, 0, 0, 0, 1, 1),
		(drawing, 4236, 4236, 0, 0, 0, 0, 1, 1),
		(drawing, 4235, 4235, 0, 0, 0, 0, 1, 1),
		(drawing, 4234, 4234, 0, 0, 0, 0, 1, 1),
		(drawing, 4233, 4233, 0, 0, 0, 0, 1, 1),
		(drawing, 4232, 4232, 0, 0, 0, 0, 1, 1),
		(drawing, 4231, 4231, 0, 0, 0, 0, 1, 1),
		(drawing, 4230, 4230, 0, 0, 0, 0, 1, 1),
		(drawing, 4229, 4229, 0, 0, 0, 0, 1, 1),
		(drawing, 4228, 4228, 0, 0, 0, 0, 1, 1),
		(drawing, 4227, 4227, 0, 0, 0, 0, 1, 1),
		(drawing, 4226, 4226, 0, 0, 0, 0, 1, 1),
		(drawing, 4225, 4225, 0, 0, 0, 0, 1, 1),
		(drawing, 4224, 4224, 0, 0, 0, 0, 1, 1),
		(drawing, 4223, 4223, 0, 0, 0, 0, 1, 1),
		(drawing, 4222, 4222, 0, 0, 0, 0, 1, 1),
		(drawing, 4221, 4221, 0, 0, 0, 0, 1, 1),
		(drawing, 4220, 4220, 0, 0, 0, 0, 1, 1),
		(drawing, 4219, 4219, 0, 0, 0, 0, 1, 1),
		(drawing, 4218, 4218, 0, 0, 0, 0, 1, 1),
		(drawing, 4217, 4217, 0, 0, 0, 0, 1, 1),
		(drawing, 4216, 4216, 0, 0, 0, 0, 1, 1),
		(drawing, 4215, 4215, 0, 0, 0, 0, 1, 1),
		(drawing, 4214, 4214, 0, 0, 0, 0, 1, 1),
		(drawing, 4213, 4213, 0, 0, 0, 0, 1, 1),
		(drawing, 4212, 4212, 0, 0, 0, 0, 1, 1),
		(drawing, 4211, 4211, 0, 0, 0, 0, 1, 1),
		(drawing, 4210, 4210, 0, 0, 0, 0, 1, 1),
		(drawing, 4209, 4209, 0, 0, 0, 0, 1, 1),
		(drawing, 4208, 4208, 0, 0, 0, 0, 1, 1),
		(drawing, 4207, 4207, 0, 0, 0, 0, 1, 1),
		(drawing, 4206, 4206, 0, 0, 0, 0, 1, 1),
		(drawing, 4205, 4205, 0, 0, 0, 0, 1, 1),
		(drawing, 4204, 4204, 0, 0, 0, 0, 1, 1),
		(drawing, 4203, 4203, 0, 0, 0, 0, 1, 1),
		(drawing, 4202, 4202, 0, 0, 0, 0, 1, 1),
		(drawing, 4201, 4201, 0, 0, 0, 0, 1, 1),
		(drawing, 4200, 4200, 0, 0, 0, 0, 1, 1),
		(drawing, 4199, 4199, 0, 0, 0, 0, 1, 1),
		(drawing, 4198, 4198, 0, 0, 0, 0, 1, 1),
		(drawing, 4197, 4197, 0, 0, 0, 0, 1, 1),
		(drawing, 4196, 4196, 0, 0, 0, 0, 1, 1),
		(drawing, 4195, 4195, 0, 0, 0, 0, 1, 1),
		(drawing, 4194, 4194, 0, 0, 0, 0, 1, 1),
		(drawing, 4193, 4193, 0, 0, 0, 0, 1, 1),
		(drawing, 4192, 4192, 0, 0, 0, 0, 1, 1),
		(drawing, 4191, 4191, 0, 0, 0, 0, 1, 1),
		(drawing, 4190, 4190, 0, 0, 0, 0, 1, 1),
		(drawing, 4189, 4189, 0, 0, 0, 0, 1, 1),
		(drawing, 4188, 4188, 0, 0, 0, 0, 1, 1),
		(drawing, 4187, 4187, 0, 0, 0, 0, 1, 1),
		(drawing, 4186, 4186, 0, 0, 0, 0, 1, 1),
		(drawing, 4185, 4185, 0, 0, 0, 0, 1, 1),
		(drawing, 4184, 4184, 0, 0, 0, 0, 1, 1),
		(drawing, 4183, 4183, 0, 0, 0, 0, 1, 1),
		(drawing, 4182, 4182, 0, 0, 0, 0, 1, 1),
		(drawing, 4181, 4181, 0, 0, 0, 0, 1, 1),
		(drawing, 4180, 4180, 0, 0, 0, 0, 1, 1),
		(drawing, 4179, 4179, 0, 0, 0, 0, 1, 1),
		(drawing, 4178, 4178, 0, 0, 0, 0, 1, 1),
		(drawing, 4177, 4177, 0, 0, 0, 0, 1, 1),
		(drawing, 4176, 4176, 0, 0, 0, 0, 1, 1),
		(drawing, 4175, 4175, 0, 0, 0, 0, 1, 1),
		(drawing, 4174, 4174, 0, 0, 0, 0, 1, 1),
		(drawing, 4173, 4173, 0, 0, 0, 0, 1, 1),
		(drawing, 4172, 4172, 0, 0, 0, 0, 1, 1),
		(drawing, 4171, 4171, 0, 0, 0, 0, 1, 1),
		(drawing, 4170, 4170, 0, 0, 0, 0, 1, 1),
		(drawing, 4169, 4169, 0, 0, 0, 0, 1, 1),
		(drawing, 4168, 4168, 0, 0, 0, 0, 1, 1),
		(drawing, 4167, 4167, 0, 0, 0, 0, 1, 1),
		(drawing, 4166, 4166, 0, 0, 0, 0, 1, 1),
		(drawing, 4165, 4165, 0, 0, 0, 0, 1, 1),
		(drawing, 4164, 4164, 0, 0, 0, 0, 1, 1),
		(drawing, 4163, 4163, 0, 0, 0, 0, 1, 1),
		(drawing, 4162, 4162, 0, 0, 0, 0, 1, 1),
		(drawing, 4161, 4161, 0, 0, 0, 0, 1, 1),
		(drawing, 4160, 4160, 0, 0, 0, 0, 1, 1),
		(drawing, 4159, 4159, 0, 0, 0, 0, 1, 1),
		(drawing, 4158, 4158, 0, 0, 0, 0, 1, 1),
		(drawing, 4157, 4157, 0, 0, 0, 0, 1, 1),
		(drawing, 4156, 4156, 0, 0, 0, 0, 1, 1),
		(drawing, 4155, 4155, 0, 0, 0, 0, 1, 1),
		(drawing, 4154, 4154, 0, 0, 0, 0, 1, 1),
		(drawing, 4153, 4153, 0, 0, 0, 0, 1, 1),
		(drawing, 4152, 4152, 0, 0, 0, 0, 1, 1),
		(drawing, 4151, 4151, 0, 0, 0, 0, 1, 1),
		(drawing, 4150, 4150, 0, 0, 0, 0, 1, 1),
		(drawing, 4149, 4149, 0, 0, 0, 0, 1, 1),
		(drawing, 4148, 4148, 0, 0, 0, 0, 1, 1),
		(drawing, 4147, 4147, 0, 0, 0, 0, 1, 1),
		(drawing, 4146, 4146, 0, 0, 0, 0, 1, 1),
		(drawing, 4145, 4145, 0, 0, 0, 0, 1, 1),
		(drawing, 4144, 4144, 0, 0, 0, 0, 1, 1),
		(drawing, 4143, 4143, 0, 0, 0, 0, 1, 1),
		(drawing, 4142, 4142, 0, 0, 0, 0, 1, 1),
		(drawing, 4141, 4141, 0, 0, 0, 0, 1, 1),
		(drawing, 4140, 4140, 0, 0, 0, 0, 1, 1),
		(drawing, 4139, 4139, 0, 0, 0, 0, 1, 1),
		(drawing, 4138, 4138, 0, 0, 0, 0, 1, 1),
		(drawing, 4137, 4137, 0, 0, 0, 0, 1, 1),
		(drawing, 4136, 4136, 0, 0, 0, 0, 1, 1),
		(drawing, 4135, 4135, 0, 0, 0, 0, 1, 1),
		(drawing, 4134, 4134, 0, 0, 0, 0, 1, 1),
		(drawing, 4133, 4133, 0, 0, 0, 0, 1, 1),
		(drawing, 4132, 4132, 0, 0, 0, 0, 1, 1),
		(drawing, 4131, 4131, 0, 0, 0, 0, 1, 1),
		(drawing, 4130, 4130, 0, 0, 0, 0, 1, 1),
		(drawing, 4129, 4129, 0, 0, 0, 0, 1, 1),
		(drawing, 4128, 4128, 0, 0, 0, 0, 1, 1),
		(drawing, 4127, 4127, 0, 0, 0, 0, 1, 1),
		(drawing, 4126, 4126, 0, 0, 0, 0, 1, 1),
		(drawing, 4125, 4125, 0, 0, 0, 0, 1, 1),
		(drawing, 4124, 4124, 0, 0, 0, 0, 1, 1),
		(drawing, 4123, 4123, 0, 0, 0, 0, 1, 1),
		(drawing, 4122, 4122, 0, 0, 0, 0, 1, 1),
		(drawing, 4121, 4121, 0, 0, 0, 0, 1, 1),
		(drawing, 4120, 4120, 0, 0, 0, 0, 1, 1),
		(drawing, 4119, 4119, 0, 0, 0, 0, 1, 1),
		(drawing, 4118, 4118, 0, 0, 0, 0, 1, 1),
		(drawing, 4117, 4117, 0, 0, 0, 0, 1, 1),
		(drawing, 4116, 4116, 0, 0, 0, 0, 1, 1),
		(drawing, 4115, 4115, 0, 0, 0, 0, 1, 1),
		(drawing, 4114, 4114, 0, 0, 0, 0, 1, 1),
		(drawing, 4113, 4113, 0, 0, 0, 0, 1, 1),
		(drawing, 4112, 4112, 0, 0, 0, 0, 1, 1),
		(drawing, 4111, 4111, 0, 0, 0, 0, 1, 1),
		(drawing, 4110, 4110, 0, 0, 0, 0, 1, 1),
		(drawing, 4109, 4109, 0, 0, 0, 0, 1, 1),
		(drawing, 4108, 4108, 0, 0, 0, 0, 1, 1),
		(drawing, 4107, 4107, 0, 0, 0, 0, 1, 1),
		(drawing, 4106, 4106, 0, 0, 0, 0, 1, 1),
		(drawing, 4105, 4105, 0, 0, 0, 0, 1, 1),
		(drawing, 4104, 4104, 0, 0, 0, 0, 1, 1),
		(drawing, 4103, 4103, 0, 0, 0, 0, 1, 1),
		(drawing, 4102, 4102, 0, 0, 0, 0, 1, 1),
		(drawing, 4101, 4101, 0, 0, 0, 0, 1, 1),
		(drawing, 4100, 4100, 0, 0, 0, 0, 1, 1),
		(drawing, 4099, 4099, 0, 0, 0, 0, 1, 1),
		(drawing, 4098, 4098, 0, 0, 0, 0, 1, 1),
		(drawing, 4097, 4097, 0, 0, 0, 0, 1, 1),
		(drawing, 4096, 4096, 0, 0, 0, 0, 1, 1),
		(drawing, 4095, 4095, 0, 0, 0, 0, 1, 1),
		(drawing, 4094, 4094, 0, 0, 0, 0, 1, 1),
		(drawing, 4093, 4093, 0, 0, 0, 0, 1, 1),
		(drawing, 4092, 4092, 0, 0, 0, 0, 1, 1),
		(drawing, 4091, 4091, 0, 0, 0, 0, 1, 1),
		(drawing, 4090, 4090, 0, 0, 0, 0, 1, 1),
		(drawing, 4089, 4089, 0, 0, 0, 0, 1, 1),
		(drawing, 4088, 4088, 0, 0, 0, 0, 1, 1),
		(drawing, 4087, 4087, 0, 0, 0, 0, 1, 1),
		(drawing, 4086, 4086, 0, 0, 0, 0, 1, 1),
		(drawing, 4085, 4085, 0, 0, 0, 0, 1, 1),
		(drawing, 4084, 4084, 0, 0, 0, 0, 1, 1),
		(drawing, 4083, 4083, 0, 0, 0, 0, 1, 1),
		(drawing, 4082, 4082, 0, 0, 0, 0, 1, 1),
		(drawing, 4081, 4081, 0, 0, 0, 0, 1, 1),
		(drawing, 4080, 4080, 0, 0, 0, 0, 1, 1),
		(drawing, 4079, 4079, 0, 0, 0, 0, 1, 1),
		(drawing, 4078, 4078, 0, 0, 0, 0, 1, 1),
		(drawing, 4077, 4077, 0, 0, 0, 0, 1, 1),
		(drawing, 4076, 4076, 0, 0, 0, 0, 1, 1),
		(drawing, 4075, 4075, 0, 0, 0, 0, 1, 1),
		(drawing, 4074, 4074, 0, 0, 0, 0, 1, 1),
		(drawing, 4073, 4073, 0, 0, 0, 0, 1, 1),
		(drawing, 4072, 4072, 0, 0, 0, 0, 1, 1),
		(drawing, 4071, 4071, 0, 0, 0, 0, 1, 1),
		(drawing, 4070, 4070, 0, 0, 0, 0, 1, 1),
		(drawing, 4069, 4069, 0, 0, 0, 0, 1, 1),
		(drawing, 4068, 4068, 0, 0, 0, 0, 1, 1),
		(drawing, 4067, 4067, 0, 0, 0, 0, 1, 1),
		(drawing, 4066, 4066, 0, 0, 0, 0, 1, 1),
		(drawing, 4065, 4065, 0, 0, 0, 0, 1, 1),
		(drawing, 4064, 4064, 0, 0, 0, 0, 1, 1),
		(drawing, 4063, 4063, 0, 0, 0, 0, 1, 1),
		(drawing, 4062, 4062, 0, 0, 0, 0, 1, 1),
		(drawing, 4061, 4061, 0, 0, 0, 0, 1, 1),
		(drawing, 4060, 4060, 0, 0, 0, 0, 1, 1),
		(drawing, 4059, 4059, 0, 0, 0, 0, 1, 1),
		(drawing, 4058, 4058, 0, 0, 0, 0, 1, 1),
		(drawing, 4057, 4057, 0, 0, 0, 0, 1, 1),
		(drawing, 4056, 4056, 0, 0, 0, 0, 1, 1),
		(drawing, 4055, 4055, 0, 0, 0, 0, 1, 1),
		(drawing, 4054, 4054, 0, 0, 0, 0, 1, 1),
		(drawing, 4053, 4053, 0, 0, 0, 0, 1, 1),
		(drawing, 4052, 4052, 0, 0, 0, 0, 1, 1),
		(drawing, 4051, 4051, 0, 0, 0, 0, 1, 1),
		(drawing, 4050, 4050, 0, 0, 0, 0, 1, 1),
		(drawing, 4049, 4049, 0, 0, 0, 0, 1, 1),
		(drawing, 4048, 4048, 0, 0, 0, 0, 1, 1),
		(drawing, 4047, 4047, 0, 0, 0, 0, 1, 1),
		(drawing, 4046, 4046, 0, 0, 0, 0, 1, 1),
		(drawing, 4045, 4045, 0, 0, 0, 0, 1, 1),
		(drawing, 4044, 4044, 0, 0, 0, 0, 1, 1),
		(drawing, 4043, 4043, 0, 0, 0, 0, 1, 1),
		(drawing, 4042, 4042, 0, 0, 0, 0, 1, 1),
		(drawing, 4041, 4041, 0, 0, 0, 0, 1, 1),
		(drawing, 4040, 4040, 0, 0, 0, 0, 1, 1),
		(drawing, 4039, 4039, 0, 0, 0, 0, 1, 1),
		(drawing, 4038, 4038, 0, 0, 0, 0, 1, 1),
		(drawing, 4037, 4037, 0, 0, 0, 0, 1, 1),
		(drawing, 4036, 4036, 0, 0, 0, 0, 1, 1),
		(drawing, 4035, 4035, 0, 0, 0, 0, 1, 1),
		(drawing, 4034, 4034, 0, 0, 0, 0, 1, 1),
		(drawing, 4033, 4033, 0, 0, 0, 0, 1, 1),
		(drawing, 4032, 4032, 0, 0, 0, 0, 1, 1),
		(drawing, 4031, 4031, 0, 0, 0, 0, 1, 1),
		(drawing, 4030, 4030, 0, 0, 0, 0, 1, 1),
		(drawing, 4029, 4029, 0, 0, 0, 0, 1, 1),
		(drawing, 4028, 4028, 0, 0, 0, 0, 1, 1),
		(drawing, 4027, 4027, 0, 0, 0, 0, 1, 1),
		(drawing, 4026, 4026, 0, 0, 0, 0, 1, 1),
		(drawing, 4025, 4025, 0, 0, 0, 0, 1, 1),
		(drawing, 4024, 4024, 0, 0, 0, 0, 1, 1),
		(drawing, 4023, 4023, 0, 0, 0, 0, 1, 1),
		(drawing, 4022, 4022, 0, 0, 0, 0, 1, 1),
		(drawing, 4021, 4021, 0, 0, 0, 0, 1, 1),
		(drawing, 4020, 4020, 0, 0, 0, 0, 1, 1),
		(drawing, 4019, 4019, 0, 0, 0, 0, 1, 1),
		(drawing, 4018, 4018, 0, 0, 0, 0, 1, 1),
		(drawing, 4017, 4017, 0, 0, 0, 0, 1, 1),
		(drawing, 4016, 4016, 0, 0, 0, 0, 1, 1),
		(drawing, 4015, 4015, 0, 0, 0, 0, 1, 1),
		(drawing, 4014, 4014, 0, 0, 0, 0, 1, 1),
		(drawing, 4013, 4013, 0, 0, 0, 0, 1, 1),
		(drawing, 4012, 4012, 0, 0, 0, 0, 1, 1),
		(drawing, 4011, 4011, 0, 0, 0, 0, 1, 1),
		(drawing, 4010, 4010, 0, 0, 0, 0, 1, 1),
		(drawing, 4009, 4009, 0, 0, 0, 0, 1, 1),
		(drawing, 4008, 4008, 0, 0, 0, 0, 1, 1),
		(drawing, 4007, 4007, 0, 0, 0, 0, 1, 1),
		(drawing, 4006, 4006, 0, 0, 0, 0, 1, 1),
		(drawing, 4005, 4005, 0, 0, 0, 0, 1, 1),
		(drawing, 4004, 4004, 0, 0, 0, 0, 1, 1),
		(drawing, 4003, 4003, 0, 0, 0, 0, 1, 1),
		(drawing, 4002, 4002, 0, 0, 0, 0, 1, 1),
		(drawing, 4001, 4001, 0, 0, 0, 0, 1, 1),
		(drawing, 4000, 4000, 0, 0, 0, 0, 1, 1),
		(drawing, 3999, 3999, 0, 0, 0, 0, 1, 1),
		(drawing, 3998, 3998, 0, 0, 0, 0, 1, 1),
		(drawing, 3997, 3997, 0, 0, 0, 0, 1, 1),
		(drawing, 3996, 3996, 0, 0, 0, 0, 1, 1),
		(drawing, 3995, 3995, 0, 0, 0, 0, 1, 1),
		(drawing, 3994, 3994, 0, 0, 0, 0, 1, 1),
		(drawing, 3993, 3993, 0, 0, 0, 0, 1, 1),
		(drawing, 3992, 3992, 0, 0, 0, 0, 1, 1),
		(drawing, 3991, 3991, 0, 0, 0, 0, 1, 1),
		(drawing, 3990, 3990, 0, 0, 0, 0, 1, 1),
		(drawing, 3989, 3989, 0, 0, 0, 0, 1, 1),
		(drawing, 3988, 3988, 0, 0, 0, 0, 1, 1),
		(drawing, 3987, 3987, 0, 0, 0, 0, 1, 1),
		(drawing, 3986, 3986, 0, 0, 0, 0, 1, 1),
		(drawing, 3985, 3985, 0, 0, 0, 0, 1, 1),
		(drawing, 3984, 3984, 0, 0, 0, 0, 1, 1),
		(drawing, 3983, 3983, 0, 0, 0, 0, 1, 1),
		(drawing, 3982, 3982, 0, 0, 0, 0, 1, 1),
		(drawing, 3981, 3981, 0, 0, 0, 0, 1, 1),
		(drawing, 3980, 3980, 0, 0, 0, 0, 1, 1),
		(drawing, 3979, 3979, 0, 0, 0, 0, 1, 1),
		(drawing, 3978, 3978, 0, 0, 0, 0, 1, 1),
		(drawing, 3977, 3977, 0, 0, 0, 0, 1, 1),
		(drawing, 3976, 3976, 0, 0, 0, 0, 1, 1),
		(drawing, 3975, 3975, 0, 0, 0, 0, 1, 1),
		(drawing, 3974, 3974, 0, 0, 0, 0, 1, 1),
		(drawing, 3973, 3973, 0, 0, 0, 0, 1, 1),
		(drawing, 3972, 3972, 0, 0, 0, 0, 1, 1),
		(drawing, 3971, 3971, 0, 0, 0, 0, 1, 1),
		(drawing, 3970, 3970, 0, 0, 0, 0, 1, 1),
		(drawing, 3969, 3969, 0, 0, 0, 0, 1, 1),
		(drawing, 3968, 3968, 0, 0, 0, 0, 1, 1),
		(drawing, 3967, 3967, 0, 0, 0, 0, 1, 1),
		(drawing, 3966, 3966, 0, 0, 0, 0, 1, 1),
		(drawing, 3965, 3965, 0, 0, 0, 0, 1, 1),
		(drawing, 3964, 3964, 0, 0, 0, 0, 1, 1),
		(drawing, 3963, 3963, 0, 0, 0, 0, 1, 1),
		(drawing, 3962, 3962, 0, 0, 0, 0, 1, 1),
		(drawing, 3961, 3961, 0, 0, 0, 0, 1, 1),
		(drawing, 3960, 3960, 0, 0, 0, 0, 1, 1),
		(drawing, 3959, 3959, 0, 0, 0, 0, 1, 1),
		(drawing, 3958, 3958, 0, 0, 0, 0, 1, 1),
		(drawing, 3957, 3957, 0, 0, 0, 0, 1, 1),
		(drawing, 3956, 3956, 0, 0, 0, 0, 1, 1),
		(drawing, 3955, 3955, 0, 0, 0, 0, 1, 1),
		(drawing, 3954, 3954, 0, 0, 0, 0, 1, 1),
		(drawing, 3953, 3953, 0, 0, 0, 0, 1, 1),
		(drawing, 3952, 3952, 0, 0, 0, 0, 1, 1),
		(drawing, 3951, 3951, 0, 0, 0, 0, 1, 1),
		(drawing, 3950, 3950, 0, 0, 0, 0, 1, 1),
		(drawing, 3949, 3949, 0, 0, 0, 0, 1, 1),
		(drawing, 3948, 3948, 0, 0, 0, 0, 1, 1),
		(drawing, 3947, 3947, 0, 0, 0, 0, 1, 1),
		(drawing, 3946, 3946, 0, 0, 0, 0, 1, 1),
		(drawing, 3945, 3945, 0, 0, 0, 0, 1, 1),
		(drawing, 3944, 3944, 0, 0, 0, 0, 1, 1),
		(drawing, 3943, 3943, 0, 0, 0, 0, 1, 1),
		(drawing, 3942, 3942, 0, 0, 0, 0, 1, 1),
		(drawing, 3941, 3941, 0, 0, 0, 0, 1, 1),
		(drawing, 3940, 3940, 0, 0, 0, 0, 1, 1),
		(drawing, 3939, 3939, 0, 0, 0, 0, 1, 1),
		(drawing, 3938, 3938, 0, 0, 0, 0, 1, 1),
		(drawing, 3937, 3937, 0, 0, 0, 0, 1, 1),
		(drawing, 3936, 3936, 0, 0, 0, 0, 1, 1),
		(drawing, 3935, 3935, 0, 0, 0, 0, 1, 1),
		(drawing, 3934, 3934, 0, 0, 0, 0, 1, 1),
		(drawing, 3933, 3933, 0, 0, 0, 0, 1, 1),
		(drawing, 3932, 3932, 0, 0, 0, 0, 1, 1),
		(drawing, 3931, 3931, 0, 0, 0, 0, 1, 1),
		(drawing, 3930, 3930, 0, 0, 0, 0, 1, 1),
		(drawing, 3929, 3929, 0, 0, 0, 0, 1, 1),
		(drawing, 3928, 3928, 0, 0, 0, 0, 1, 1),
		(drawing, 3927, 3927, 0, 0, 0, 0, 1, 1),
		(drawing, 3926, 3926, 0, 0, 0, 0, 1, 1),
		(drawing, 3925, 3925, 0, 0, 0, 0, 1, 1),
		(drawing, 3924, 3924, 0, 0, 0, 0, 1, 1),
		(drawing, 3923, 3923, 0, 0, 0, 0, 1, 1),
		(drawing, 3922, 3922, 0, 0, 0, 0, 1, 1),
		(drawing, 3921, 3921, 0, 0, 0, 0, 1, 1),
		(drawing, 3920, 3920, 0, 0, 0, 0, 1, 1),
		(drawing, 3919, 3919, 0, 0, 0, 0, 1, 1),
		(drawing, 3918, 3918, 0, 0, 0, 0, 1, 1),
		(drawing, 3917, 3917, 0, 0, 0, 0, 1, 1),
		(drawing, 3916, 3916, 0, 0, 0, 0, 1, 1),
		(drawing, 3915, 3915, 0, 0, 0, 0, 1, 1),
		(drawing, 3914, 3914, 0, 0, 0, 0, 1, 1),
		(drawing, 3913, 3913, 0, 0, 0, 0, 1, 1),
		(drawing, 3912, 3912, 0, 0, 0, 0, 1, 1),
		(drawing, 3911, 3911, 0, 0, 0, 0, 1, 1),
		(drawing, 3910, 3910, 0, 0, 0, 0, 1, 1),
		(drawing, 3909, 3909, 0, 0, 0, 0, 1, 1),
		(drawing, 3908, 3908, 0, 0, 0, 0, 1, 1),
		(drawing, 3907, 3907, 0, 0, 0, 0, 1, 1),
		(drawing, 3906, 3906, 0, 0, 0, 0, 1, 1),
		(drawing, 3905, 3905, 0, 0, 0, 0, 1, 1),
		(drawing, 3904, 3904, 0, 0, 0, 0, 1, 1),
		(drawing, 3903, 3903, 0, 0, 0, 0, 1, 1),
		(drawing, 3902, 3902, 0, 0, 0, 0, 1, 1),
		(drawing, 3901, 3901, 0, 0, 0, 0, 1, 1),
		(drawing, 3900, 3900, 0, 0, 0, 0, 1, 1),
		(drawing, 3899, 3899, 0, 0, 0, 0, 1, 1),
		(drawing, 3898, 3898, 0, 0, 0, 0, 1, 1),
		(drawing, 3897, 3897, 0, 0, 0, 0, 1, 1),
		(drawing, 3896, 3896, 0, 0, 0, 0, 1, 1),
		(drawing, 3895, 3895, 0, 0, 0, 0, 1, 1),
		(drawing, 3894, 3894, 0, 0, 0, 0, 1, 1),
		(drawing, 3893, 3893, 0, 0, 0, 0, 1, 1),
		(drawing, 3892, 3892, 0, 0, 0, 0, 1, 1),
		(drawing, 3891, 3891, 0, 0, 0, 0, 1, 1),
		(drawing, 3890, 3890, 0, 0, 0, 0, 1, 1),
		(drawing, 3889, 3889, 0, 0, 0, 0, 1, 1),
		(drawing, 3888, 3888, 0, 0, 0, 0, 1, 1),
		(drawing, 3887, 3887, 0, 0, 0, 0, 1, 1),
		(drawing, 3886, 3886, 0, 0, 0, 0, 1, 1),
		(drawing, 3885, 3885, 0, 0, 0, 0, 1, 1),
		(drawing, 3884, 3884, 0, 0, 0, 0, 1, 1),
		(drawing, 3883, 3883, 0, 0, 0, 0, 1, 1),
		(drawing, 3882, 3882, 0, 0, 0, 0, 1, 1),
		(drawing, 3881, 3881, 0, 0, 0, 0, 1, 1),
		(drawing, 3880, 3880, 0, 0, 0, 0, 1, 1),
		(drawing, 3879, 3879, 0, 0, 0, 0, 1, 1),
		(drawing, 3878, 3878, 0, 0, 0, 0, 1, 1),
		(drawing, 3877, 3877, 0, 0, 0, 0, 1, 1),
		(drawing, 3876, 3876, 0, 0, 0, 0, 1, 1),
		(drawing, 3875, 3875, 0, 0, 0, 0, 1, 1),
		(drawing, 3874, 3874, 0, 0, 0, 0, 1, 1),
		(drawing, 3873, 3873, 0, 0, 0, 0, 1, 1),
		(drawing, 3872, 3872, 0, 0, 0, 0, 1, 1),
		(drawing, 3871, 3871, 0, 0, 0, 0, 1, 1),
		(drawing, 3870, 3870, 0, 0, 0, 0, 1, 1),
		(drawing, 3869, 3869, 0, 0, 0, 0, 1, 1),
		(drawing, 3868, 3868, 0, 0, 0, 0, 1, 1),
		(drawing, 3867, 3867, 0, 0, 0, 0, 1, 1),
		(drawing, 3866, 3866, 0, 0, 0, 0, 1, 1),
		(drawing, 3865, 3865, 0, 0, 0, 0, 1, 1),
		(drawing, 3864, 3864, 0, 0, 0, 0, 1, 1),
		(drawing, 3863, 3863, 0, 0, 0, 0, 1, 1),
		(drawing, 3862, 3862, 0, 0, 0, 0, 1, 1),
		(drawing, 3861, 3861, 0, 0, 0, 0, 1, 1),
		(drawing, 3860, 3860, 0, 0, 0, 0, 1, 1),
		(drawing, 3859, 3859, 0, 0, 0, 0, 1, 1),
		(drawing, 3858, 3858, 0, 0, 0, 0, 1, 1),
		(drawing, 3857, 3857, 0, 0, 0, 0, 1, 1),
		(drawing, 3856, 3856, 0, 0, 0, 0, 1, 1),
		(drawing, 3855, 3855, 0, 0, 0, 0, 1, 1),
		(drawing, 3854, 3854, 0, 0, 0, 0, 1, 1),
		(drawing, 3853, 3853, 0, 0, 0, 0, 1, 1),
		(drawing, 3852, 3852, 0, 0, 0, 0, 1, 1),
		(drawing, 3851, 3851, 0, 0, 0, 0, 1, 1),
		(drawing, 3850, 3850, 0, 0, 0, 0, 1, 1),
		(drawing, 3849, 3849, 0, 0, 0, 0, 1, 1),
		(drawing, 3848, 3848, 0, 0, 0, 0, 1, 1),
		(drawing, 3847, 3847, 0, 0, 0, 0, 1, 1),
		(drawing, 3846, 3846, 0, 0, 0, 0, 1, 1),
		(drawing, 3845, 3845, 0, 0, 0, 0, 1, 1),
		(drawing, 3844, 3844, 0, 0, 0, 0, 1, 1),
		(drawing, 3843, 3843, 0, 0, 0, 0, 1, 1),
		(drawing, 3842, 3842, 0, 0, 0, 0, 1, 1),
		(drawing, 3841, 3841, 0, 0, 0, 0, 1, 1),
		(drawing, 3840, 3840, 0, 0, 0, 0, 1, 1),
		(drawing, 3839, 3839, 0, 0, 0, 0, 1, 1),
		(drawing, 3838, 3838, 0, 0, 0, 0, 1, 1),
		(drawing, 3837, 3837, 0, 0, 0, 0, 1, 1),
		(drawing, 3836, 3836, 0, 0, 0, 0, 1, 1),
		(drawing, 3835, 3835, 0, 0, 0, 0, 1, 1),
		(drawing, 3834, 3834, 0, 0, 0, 0, 1, 1),
		(drawing, 3833, 3833, 0, 0, 0, 0, 1, 1),
		(drawing, 3832, 3832, 0, 0, 0, 0, 1, 1),
		(drawing, 3831, 3831, 0, 0, 0, 0, 1, 1),
		(drawing, 3830, 3830, 0, 0, 0, 0, 1, 1),
		(drawing, 3829, 3829, 0, 0, 0, 0, 1, 1),
		(drawing, 3828, 3828, 0, 0, 0, 0, 1, 1),
		(drawing, 3827, 3827, 0, 0, 0, 0, 1, 1),
		(drawing, 3826, 3826, 0, 0, 0, 0, 1, 1),
		(drawing, 3825, 3825, 0, 0, 0, 0, 1, 1),
		(drawing, 3824, 3824, 0, 0, 0, 0, 1, 1),
		(drawing, 3823, 3823, 0, 0, 0, 0, 1, 1),
		(drawing, 3822, 3822, 0, 0, 0, 0, 1, 1),
		(drawing, 3821, 3821, 0, 0, 0, 0, 1, 1),
		(drawing, 3820, 3820, 0, 0, 0, 0, 1, 1),
		(drawing, 3819, 3819, 0, 0, 0, 0, 1, 1),
		(drawing, 3818, 3818, 0, 0, 0, 0, 1, 1),
		(drawing, 3817, 3817, 0, 0, 0, 0, 1, 1),
		(drawing, 3816, 3816, 0, 0, 0, 0, 1, 1),
		(drawing, 3815, 3815, 0, 0, 0, 0, 1, 1),
		(drawing, 3814, 3814, 0, 0, 0, 0, 1, 1),
		(drawing, 3813, 3813, 0, 0, 0, 0, 1, 1),
		(drawing, 3812, 3812, 0, 0, 0, 0, 1, 1),
		(drawing, 3811, 3811, 0, 0, 0, 0, 1, 1),
		(drawing, 3810, 3810, 0, 0, 0, 0, 1, 1),
		(drawing, 3809, 3809, 0, 0, 0, 0, 1, 1),
		(drawing, 3808, 3808, 0, 0, 0, 0, 1, 1),
		(drawing, 3807, 3807, 0, 0, 0, 0, 1, 1),
		(drawing, 3806, 3806, 0, 0, 0, 0, 1, 1),
		(drawing, 3805, 3805, 0, 0, 0, 0, 1, 1),
		(drawing, 3804, 3804, 0, 0, 0, 0, 1, 1),
		(drawing, 3803, 3803, 0, 0, 0, 0, 1, 1),
		(drawing, 3802, 3802, 0, 0, 0, 0, 1, 1),
		(drawing, 3801, 3801, 0, 0, 0, 0, 1, 1),
		(drawing, 3800, 3800, 0, 0, 0, 0, 1, 1),
		(drawing, 3799, 3799, 0, 0, 0, 0, 1, 1),
		(drawing, 3798, 3798, 0, 0, 0, 0, 1, 1),
		(drawing, 3797, 3797, 0, 0, 0, 0, 1, 1),
		(drawing, 3796, 3796, 0, 0, 0, 0, 1, 1),
		(drawing, 3795, 3795, 0, 0, 0, 0, 1, 1),
		(drawing, 3794, 3794, 0, 0, 0, 0, 1, 1),
		(drawing, 3793, 3793, 0, 0, 0, 0, 1, 1),
		(drawing, 3792, 3792, 0, 0, 0, 0, 1, 1),
		(drawing, 3791, 3791, 0, 0, 0, 0, 1, 1),
		(drawing, 3790, 3790, 0, 0, 0, 0, 1, 1),
		(drawing, 3789, 3789, 0, 0, 0, 0, 1, 1),
		(drawing, 3788, 3788, 0, 0, 0, 0, 1, 1),
		(drawing, 3787, 3787, 0, 0, 0, 0, 1, 1),
		(drawing, 3786, 3786, 0, 0, 0, 0, 1, 1),
		(drawing, 3785, 3785, 0, 0, 0, 0, 1, 1),
		(drawing, 3784, 3784, 0, 0, 0, 0, 1, 1),
		(drawing, 3783, 3783, 0, 0, 0, 0, 1, 1),
		(drawing, 3782, 3782, 0, 0, 0, 0, 1, 1),
		(drawing, 3781, 3781, 0, 0, 0, 0, 1, 1),
		(drawing, 3780, 3780, 0, 0, 0, 0, 1, 1),
		(drawing, 3779, 3779, 0, 0, 0, 0, 1, 1),
		(drawing, 3778, 3778, 0, 0, 0, 0, 1, 1),
		(drawing, 3777, 3777, 0, 0, 0, 0, 1, 1),
		(drawing, 3776, 3776, 0, 0, 0, 0, 1, 1),
		(drawing, 3775, 3775, 0, 0, 0, 0, 1, 1),
		(drawing, 3774, 3774, 0, 0, 0, 0, 1, 1),
		(drawing, 3773, 3773, 0, 0, 0, 0, 1, 1),
		(drawing, 3772, 3772, 0, 0, 0, 0, 1, 1),
		(drawing, 3771, 3771, 0, 0, 0, 0, 1, 1),
		(drawing, 3770, 3770, 0, 0, 0, 0, 1, 1),
		(drawing, 3769, 3769, 0, 0, 0, 0, 1, 1),
		(drawing, 3768, 3768, 0, 0, 0, 0, 1, 1),
		(drawing, 3767, 3767, 0, 0, 0, 0, 1, 1),
		(drawing, 3766, 3766, 0, 0, 0, 0, 1, 1),
		(drawing, 3765, 3765, 0, 0, 0, 0, 1, 1),
		(drawing, 3764, 3764, 0, 0, 0, 0, 1, 1),
		(drawing, 3763, 3763, 0, 0, 0, 0, 1, 1),
		(drawing, 3762, 3762, 0, 0, 0, 0, 1, 1),
		(drawing, 3761, 3761, 0, 0, 0, 0, 1, 1),
		(drawing, 3760, 3760, 0, 0, 0, 0, 1, 1),
		(drawing, 3759, 3759, 0, 0, 0, 0, 1, 1),
		(drawing, 3758, 3758, 0, 0, 0, 0, 1, 1),
		(drawing, 3757, 3757, 0, 0, 0, 0, 1, 1),
		(drawing, 3756, 3756, 0, 0, 0, 0, 1, 1),
		(drawing, 3755, 3755, 0, 0, 0, 0, 1, 1),
		(drawing, 3754, 3754, 0, 0, 0, 0, 1, 1),
		(drawing, 3753, 3753, 0, 0, 0, 0, 1, 1),
		(drawing, 3752, 3752, 0, 0, 0, 0, 1, 1),
		(drawing, 3751, 3751, 0, 0, 0, 0, 1, 1),
		(drawing, 3750, 3750, 0, 0, 0, 0, 1, 1),
		(drawing, 3749, 3749, 0, 0, 0, 0, 1, 1),
		(drawing, 3748, 3748, 0, 0, 0, 0, 1, 1),
		(drawing, 3747, 3747, 0, 0, 0, 0, 1, 1),
		(drawing, 3746, 3746, 0, 0, 0, 0, 1, 1),
		(drawing, 3745, 3745, 0, 0, 0, 0, 1, 1),
		(drawing, 3744, 3744, 0, 0, 0, 0, 1, 1),
		(drawing, 3743, 3743, 0, 0, 0, 0, 1, 1),
		(drawing, 3742, 3742, 0, 0, 0, 0, 1, 1),
		(drawing, 3741, 3741, 0, 0, 0, 0, 1, 1),
		(drawing, 3740, 3740, 0, 0, 0, 0, 1, 1),
		(drawing, 3739, 3739, 0, 0, 0, 0, 1, 1),
		(drawing, 3738, 3738, 0, 0, 0, 0, 1, 1),
		(drawing, 3737, 3737, 0, 0, 0, 0, 1, 1),
		(drawing, 3736, 3736, 0, 0, 0, 0, 1, 1),
		(drawing, 3735, 3735, 0, 0, 0, 0, 1, 1),
		(drawing, 3734, 3734, 0, 0, 0, 0, 1, 1),
		(drawing, 3733, 3733, 0, 0, 0, 0, 1, 1),
		(drawing, 3732, 3732, 0, 0, 0, 0, 1, 1),
		(drawing, 3731, 3731, 0, 0, 0, 0, 1, 1),
		(drawing, 3730, 3730, 0, 0, 0, 0, 1, 1),
		(drawing, 3729, 3729, 0, 0, 0, 0, 1, 1),
		(drawing, 3728, 3728, 0, 0, 0, 0, 1, 1),
		(drawing, 3727, 3727, 0, 0, 0, 0, 1, 1),
		(drawing, 3726, 3726, 0, 0, 0, 0, 1, 1),
		(drawing, 3725, 3725, 0, 0, 0, 0, 1, 1),
		(drawing, 3724, 3724, 0, 0, 0, 0, 1, 1),
		(drawing, 3723, 3723, 0, 0, 0, 0, 1, 1),
		(drawing, 3722, 3722, 0, 0, 0, 0, 1, 1),
		(drawing, 3721, 3721, 0, 0, 0, 0, 1, 1),
		(drawing, 3720, 3720, 0, 0, 0, 0, 1, 1),
		(drawing, 3719, 3719, 0, 0, 0, 0, 1, 1),
		(drawing, 3718, 3718, 0, 0, 0, 0, 1, 1),
		(drawing, 3717, 3717, 0, 0, 0, 0, 1, 1),
		(drawing, 3716, 3716, 0, 0, 0, 0, 1, 1),
		(drawing, 3715, 3715, 0, 0, 0, 0, 1, 1),
		(drawing, 3714, 3714, 0, 0, 0, 0, 1, 1),
		(drawing, 3713, 3713, 0, 0, 0, 0, 1, 1),
		(drawing, 3712, 3712, 0, 0, 0, 0, 1, 1),
		(drawing, 3711, 3711, 0, 0, 0, 0, 1, 1),
		(drawing, 3710, 3710, 0, 0, 0, 0, 1, 1),
		(drawing, 3709, 3709, 0, 0, 0, 0, 1, 1),
		(drawing, 3708, 3708, 0, 0, 0, 0, 1, 1),
		(drawing, 3707, 3707, 0, 0, 0, 0, 1, 1),
		(drawing, 3706, 3706, 0, 0, 0, 0, 1, 1),
		(drawing, 3705, 3705, 0, 0, 0, 0, 1, 1),
		(drawing, 3704, 3704, 0, 0, 0, 0, 1, 1),
		(drawing, 3703, 3703, 0, 0, 0, 0, 1, 1),
		(drawing, 3702, 3702, 0, 0, 0, 0, 1, 1),
		(drawing, 3701, 3701, 0, 0, 0, 0, 1, 1),
		(drawing, 3700, 3700, 0, 0, 0, 0, 1, 1),
		(drawing, 3699, 3699, 0, 0, 0, 0, 1, 1),
		(drawing, 3698, 3698, 0, 0, 0, 0, 1, 1),
		(drawing, 3697, 3697, 0, 0, 0, 0, 1, 1),
		(drawing, 3696, 3696, 0, 0, 0, 0, 1, 1),
		(drawing, 3695, 3695, 0, 0, 0, 0, 1, 1),
		(drawing, 3694, 3694, 0, 0, 0, 0, 1, 1),
		(drawing, 3693, 3693, 0, 0, 0, 0, 1, 1),
		(drawing, 3692, 3692, 0, 0, 0, 0, 1, 1),
		(drawing, 3691, 3691, 0, 0, 0, 0, 1, 1),
		(drawing, 3690, 3690, 0, 0, 0, 0, 1, 1),
		(drawing, 3689, 3689, 0, 0, 0, 0, 1, 1),
		(drawing, 3688, 3688, 0, 0, 0, 0, 1, 1),
		(drawing, 3687, 3687, 0, 0, 0, 0, 1, 1),
		(drawing, 3686, 3686, 0, 0, 0, 0, 1, 1),
		(drawing, 3685, 3685, 0, 0, 0, 0, 1, 1),
		(drawing, 3684, 3684, 0, 0, 0, 0, 1, 1),
		(drawing, 3683, 3683, 0, 0, 0, 0, 1, 1),
		(drawing, 3682, 3682, 0, 0, 0, 0, 1, 1),
		(drawing, 3681, 3681, 0, 0, 0, 0, 1, 1),
		(drawing, 3680, 3680, 0, 0, 0, 0, 1, 1),
		(drawing, 3679, 3679, 0, 0, 0, 0, 1, 1),
		(drawing, 3678, 3678, 0, 0, 0, 0, 1, 1),
		(drawing, 3677, 3677, 0, 0, 0, 0, 1, 1),
		(drawing, 3676, 3676, 0, 0, 0, 0, 1, 1),
		(drawing, 3675, 3675, 0, 0, 0, 0, 1, 1),
		(drawing, 3674, 3674, 0, 0, 0, 0, 1, 1),
		(drawing, 3673, 3673, 0, 0, 0, 0, 1, 1),
		(drawing, 3672, 3672, 0, 0, 0, 0, 1, 1),
		(drawing, 3671, 3671, 0, 0, 0, 0, 1, 1),
		(drawing, 3670, 3670, 0, 0, 0, 0, 1, 1),
		(drawing, 3669, 3669, 0, 0, 0, 0, 1, 1),
		(drawing, 3668, 3668, 0, 0, 0, 0, 1, 1),
		(drawing, 3667, 3667, 0, 0, 0, 0, 1, 1),
		(drawing, 3666, 3666, 0, 0, 0, 0, 1, 1),
		(drawing, 3665, 3665, 0, 0, 0, 0, 1, 1),
		(drawing, 3664, 3664, 0, 0, 0, 0, 1, 1),
		(drawing, 3663, 3663, 0, 0, 0, 0, 1, 1),
		(drawing, 3662, 3662, 0, 0, 0, 0, 1, 1),
		(drawing, 3661, 3661, 0, 0, 0, 0, 1, 1),
		(drawing, 3660, 3660, 0, 0, 0, 0, 1, 1),
		(drawing, 3659, 3659, 0, 0, 0, 0, 1, 1),
		(drawing, 3658, 3658, 0, 0, 0, 0, 1, 1),
		(drawing, 3657, 3657, 0, 0, 0, 0, 1, 1),
		(drawing, 3656, 3656, 0, 0, 0, 0, 1, 1),
		(drawing, 3655, 3655, 0, 0, 0, 0, 1, 1),
		(drawing, 3654, 3654, 0, 0, 0, 0, 1, 1),
		(drawing, 3653, 3653, 0, 0, 0, 0, 1, 1),
		(drawing, 3652, 3652, 0, 0, 0, 0, 1, 1),
		(drawing, 3651, 3651, 0, 0, 0, 0, 1, 1),
		(drawing, 3650, 3650, 0, 0, 0, 0, 1, 1),
		(drawing, 3649, 3649, 0, 0, 0, 0, 1, 1),
		(drawing, 3648, 3648, 0, 0, 0, 0, 1, 1),
		(drawing, 3647, 3647, 0, 0, 0, 0, 1, 1),
		(drawing, 3646, 3646, 0, 0, 0, 0, 1, 1),
		(drawing, 3645, 3645, 0, 0, 0, 0, 1, 1),
		(drawing, 3644, 3644, 0, 0, 0, 0, 1, 1),
		(drawing, 3643, 3643, 0, 0, 0, 0, 1, 1),
		(drawing, 3642, 3642, 0, 0, 0, 0, 1, 1),
		(drawing, 3641, 3641, 0, 0, 0, 0, 1, 1),
		(drawing, 3640, 3640, 0, 0, 0, 0, 1, 1),
		(drawing, 3639, 3639, 0, 0, 0, 0, 1, 1),
		(drawing, 3638, 3638, 0, 0, 0, 0, 1, 1),
		(drawing, 3637, 3637, 0, 0, 0, 0, 1, 1),
		(drawing, 3636, 3636, 0, 0, 0, 0, 1, 1),
		(drawing, 3635, 3635, 0, 0, 0, 0, 1, 1),
		(drawing, 3634, 3634, 0, 0, 0, 0, 1, 1),
		(drawing, 3633, 3633, 0, 0, 0, 0, 1, 1),
		(drawing, 3632, 3632, 0, 0, 0, 0, 1, 1),
		(drawing, 3631, 3631, 0, 0, 0, 0, 1, 1),
		(drawing, 3630, 3630, 0, 0, 0, 0, 1, 1),
		(drawing, 3629, 3629, 0, 0, 0, 0, 1, 1),
		(drawing, 3628, 3628, 0, 0, 0, 0, 1, 1),
		(drawing, 3627, 3627, 0, 0, 0, 0, 1, 1),
		(drawing, 3626, 3626, 0, 0, 0, 0, 1, 1),
		(drawing, 3625, 3625, 0, 0, 0, 0, 1, 1),
		(drawing, 3624, 3624, 0, 0, 0, 0, 1, 1),
		(drawing, 3623, 3623, 0, 0, 0, 0, 1, 1),
		(drawing, 3622, 3622, 0, 0, 0, 0, 1, 1),
		(drawing, 3621, 3621, 0, 0, 0, 0, 1, 1),
		(drawing, 3620, 3620, 0, 0, 0, 0, 1, 1),
		(drawing, 3619, 3619, 0, 0, 0, 0, 1, 1),
		(drawing, 3618, 3618, 0, 0, 0, 0, 1, 1),
		(drawing, 3617, 3617, 0, 0, 0, 0, 1, 1),
		(drawing, 3616, 3616, 0, 0, 0, 0, 1, 1),
		(drawing, 3615, 3615, 0, 0, 0, 0, 1, 1),
		(drawing, 3614, 3614, 0, 0, 0, 0, 1, 1),
		(drawing, 3613, 3613, 0, 0, 0, 0, 1, 1),
		(drawing, 3612, 3612, 0, 0, 0, 0, 1, 1),
		(drawing, 3611, 3611, 0, 0, 0, 0, 1, 1),
		(drawing, 3610, 3610, 0, 0, 0, 0, 1, 1),
		(drawing, 3609, 3609, 0, 0, 0, 0, 1, 1),
		(drawing, 3608, 3608, 0, 0, 0, 0, 1, 1),
		(drawing, 3607, 3607, 0, 0, 0, 0, 1, 1),
		(drawing, 3606, 3606, 0, 0, 0, 0, 1, 1),
		(drawing, 3605, 3605, 0, 0, 0, 0, 1, 1),
		(drawing, 3604, 3604, 0, 0, 0, 0, 1, 1),
		(drawing, 3603, 3603, 0, 0, 0, 0, 1, 1),
		(drawing, 3602, 3602, 0, 0, 0, 0, 1, 1),
		(drawing, 3601, 3601, 0, 0, 0, 0, 1, 1),
		(drawing, 3600, 3600, 0, 0, 0, 0, 1, 1),
		(drawing, 3599, 3599, 0, 0, 0, 0, 1, 1),
		(drawing, 3598, 3598, 0, 0, 0, 0, 1, 1),
		(drawing, 3597, 3597, 0, 0, 0, 0, 1, 1),
		(drawing, 3596, 3596, 0, 0, 0, 0, 1, 1),
		(drawing, 3595, 3595, 0, 0, 0, 0, 1, 1),
		(drawing, 3594, 3594, 0, 0, 0, 0, 1, 1),
		(drawing, 3593, 3593, 0, 0, 0, 0, 1, 1),
		(drawing, 3592, 3592, 0, 0, 0, 0, 1, 1),
		(drawing, 3591, 3591, 0, 0, 0, 0, 1, 1),
		(drawing, 3590, 3590, 0, 0, 0, 0, 1, 1),
		(drawing, 3589, 3589, 0, 0, 0, 0, 1, 1),
		(drawing, 3588, 3588, 0, 0, 0, 0, 1, 1),
		(drawing, 3587, 3587, 0, 0, 0, 0, 1, 1),
		(drawing, 3586, 3586, 0, 0, 0, 0, 1, 1),
		(drawing, 3585, 3585, 0, 0, 0, 0, 1, 1),
		(drawing, 3584, 3584, 0, 0, 0, 0, 1, 1),
		(drawing, 3583, 3583, 0, 0, 0, 0, 1, 1),
		(drawing, 3582, 3582, 0, 0, 0, 0, 1, 1),
		(drawing, 3581, 3581, 0, 0, 0, 0, 1, 1),
		(drawing, 3580, 3580, 0, 0, 0, 0, 1, 1),
		(drawing, 3579, 3579, 0, 0, 0, 0, 1, 1),
		(drawing, 3578, 3578, 0, 0, 0, 0, 1, 1),
		(drawing, 3577, 3577, 0, 0, 0, 0, 1, 1),
		(drawing, 3576, 3576, 0, 0, 0, 0, 1, 1),
		(drawing, 3575, 3575, 0, 0, 0, 0, 1, 1),
		(drawing, 3574, 3574, 0, 0, 0, 0, 1, 1),
		(drawing, 3573, 3573, 0, 0, 0, 0, 1, 1),
		(drawing, 3572, 3572, 0, 0, 0, 0, 1, 1),
		(drawing, 3571, 3571, 0, 0, 0, 0, 1, 1),
		(drawing, 3570, 3570, 0, 0, 0, 0, 1, 1),
		(drawing, 3569, 3569, 0, 0, 0, 0, 1, 1),
		(drawing, 3568, 3568, 0, 0, 0, 0, 1, 1),
		(drawing, 3567, 3567, 0, 0, 0, 0, 1, 1),
		(drawing, 3566, 3566, 0, 0, 0, 0, 1, 1),
		(drawing, 3565, 3565, 0, 0, 0, 0, 1, 1),
		(drawing, 3564, 3564, 0, 0, 0, 0, 1, 1),
		(drawing, 3563, 3563, 0, 0, 0, 0, 1, 1),
		(drawing, 3562, 3562, 0, 0, 0, 0, 1, 1),
		(drawing, 3561, 3561, 0, 0, 0, 0, 1, 1),
		(drawing, 3560, 3560, 0, 0, 0, 0, 1, 1),
		(drawing, 3559, 3559, 0, 0, 0, 0, 1, 1),
		(drawing, 3558, 3558, 0, 0, 0, 0, 1, 1),
		(drawing, 3557, 3557, 0, 0, 0, 0, 1, 1),
		(drawing, 3556, 3556, 0, 0, 0, 0, 1, 1),
		(drawing, 3555, 3555, 0, 0, 0, 0, 1, 1),
		(drawing, 3554, 3554, 0, 0, 0, 0, 1, 1),
		(drawing, 3553, 3553, 0, 0, 0, 0, 1, 1),
		(drawing, 3552, 3552, 0, 0, 0, 0, 1, 1),
		(drawing, 3551, 3551, 0, 0, 0, 0, 1, 1),
		(drawing, 3550, 3550, 0, 0, 0, 0, 1, 1),
		(drawing, 3549, 3549, 0, 0, 0, 0, 1, 1),
		(drawing, 3548, 3548, 0, 0, 0, 0, 1, 1),
		(drawing, 3547, 3547, 0, 0, 0, 0, 1, 1),
		(drawing, 3546, 3546, 0, 0, 0, 0, 1, 1),
		(drawing, 3545, 3545, 0, 0, 0, 0, 1, 1),
		(drawing, 3544, 3544, 0, 0, 0, 0, 1, 1),
		(drawing, 3543, 3543, 0, 0, 0, 0, 1, 1),
		(drawing, 3542, 3542, 0, 0, 0, 0, 1, 1),
		(drawing, 3541, 3541, 0, 0, 0, 0, 1, 1),
		(drawing, 3540, 3540, 0, 0, 0, 0, 1, 1),
		(drawing, 3539, 3539, 0, 0, 0, 0, 1, 1),
		(drawing, 3538, 3538, 0, 0, 0, 0, 1, 1),
		(drawing, 3537, 3537, 0, 0, 0, 0, 1, 1),
		(drawing, 3536, 3536, 0, 0, 0, 0, 1, 1),
		(drawing, 3535, 3535, 0, 0, 0, 0, 1, 1),
		(drawing, 3534, 3534, 0, 0, 0, 0, 1, 1),
		(drawing, 3533, 3533, 0, 0, 0, 0, 1, 1),
		(drawing, 3532, 3532, 0, 0, 0, 0, 1, 1),
		(drawing, 3531, 3531, 0, 0, 0, 0, 1, 1),
		(drawing, 3530, 3530, 0, 0, 0, 0, 1, 1),
		(drawing, 3529, 3529, 0, 0, 0, 0, 1, 1),
		(drawing, 3528, 3528, 0, 0, 0, 0, 1, 1),
		(drawing, 3527, 3527, 0, 0, 0, 0, 1, 1),
		(drawing, 3526, 3526, 0, 0, 0, 0, 1, 1),
		(drawing, 3525, 3525, 0, 0, 0, 0, 1, 1),
		(drawing, 3524, 3524, 0, 0, 0, 0, 1, 1),
		(drawing, 3523, 3523, 0, 0, 0, 0, 1, 1),
		(drawing, 3522, 3522, 0, 0, 0, 0, 1, 1),
		(drawing, 3521, 3521, 0, 0, 0, 0, 1, 1),
		(drawing, 3520, 3520, 0, 0, 0, 0, 1, 1),
		(drawing, 3519, 3519, 0, 0, 0, 0, 1, 1),
		(drawing, 3518, 3518, 0, 0, 0, 0, 1, 1),
		(drawing, 3517, 3517, 0, 0, 0, 0, 1, 1),
		(drawing, 3516, 3516, 0, 0, 0, 0, 1, 1),
		(drawing, 3515, 3515, 0, 0, 0, 0, 1, 1),
		(drawing, 3514, 3514, 0, 0, 0, 0, 1, 1),
		(drawing, 3513, 3513, 0, 0, 0, 0, 1, 1),
		(drawing, 3512, 3512, 0, 0, 0, 0, 1, 1),
		(drawing, 3511, 3511, 0, 0, 0, 0, 1, 1),
		(drawing, 3510, 3510, 0, 0, 0, 0, 1, 1),
		(drawing, 3509, 3509, 0, 0, 0, 0, 1, 1),
		(drawing, 3508, 3508, 0, 0, 0, 0, 1, 1),
		(drawing, 3507, 3507, 0, 0, 0, 0, 1, 1),
		(drawing, 3506, 3506, 0, 0, 0, 0, 1, 1),
		(drawing, 3505, 3505, 0, 0, 0, 0, 1, 1),
		(drawing, 3504, 3504, 0, 0, 0, 0, 1, 1),
		(drawing, 3503, 3503, 0, 0, 0, 0, 1, 1),
		(drawing, 3502, 3502, 0, 0, 0, 0, 1, 1),
		(drawing, 3501, 3501, 0, 0, 0, 0, 1, 1),
		(drawing, 3500, 3500, 0, 0, 0, 0, 1, 1),
		(drawing, 3499, 3499, 0, 0, 0, 0, 1, 1),
		(drawing, 3498, 3498, 0, 0, 0, 0, 1, 1),
		(drawing, 3497, 3497, 0, 0, 0, 0, 1, 1),
		(drawing, 3496, 3496, 0, 0, 0, 0, 1, 1),
		(drawing, 3495, 3495, 0, 0, 0, 0, 1, 1),
		(drawing, 3494, 3494, 0, 0, 0, 0, 1, 1),
		(drawing, 3493, 3493, 0, 0, 0, 0, 1, 1),
		(drawing, 3492, 3492, 0, 0, 0, 0, 1, 1),
		(drawing, 3491, 3491, 0, 0, 0, 0, 1, 1),
		(drawing, 3490, 3490, 0, 0, 0, 0, 1, 1),
		(drawing, 3489, 3489, 0, 0, 0, 0, 1, 1),
		(drawing, 3488, 3488, 0, 0, 0, 0, 1, 1),
		(drawing, 3487, 3487, 0, 0, 0, 0, 1, 1),
		(drawing, 3486, 3486, 0, 0, 0, 0, 1, 1),
		(drawing, 3485, 3485, 0, 0, 0, 0, 1, 1),
		(drawing, 3484, 3484, 0, 0, 0, 0, 1, 1),
		(drawing, 3483, 3483, 0, 0, 0, 0, 1, 1),
		(drawing, 3482, 3482, 0, 0, 0, 0, 1, 1),
		(drawing, 3481, 3481, 0, 0, 0, 0, 1, 1),
		(drawing, 3480, 3480, 0, 0, 0, 0, 1, 1),
		(drawing, 3479, 3479, 0, 0, 0, 0, 1, 1),
		(drawing, 3478, 3478, 0, 0, 0, 0, 1, 1),
		(drawing, 3477, 3477, 0, 0, 0, 0, 1, 1),
		(drawing, 3476, 3476, 0, 0, 0, 0, 1, 1),
		(drawing, 3475, 3475, 0, 0, 0, 0, 1, 1),
		(drawing, 3474, 3474, 0, 0, 0, 0, 1, 1),
		(drawing, 3473, 3473, 0, 0, 0, 0, 1, 1),
		(drawing, 3472, 3472, 0, 0, 0, 0, 1, 1),
		(drawing, 3471, 3471, 0, 0, 0, 0, 1, 1),
		(drawing, 3470, 3470, 0, 0, 0, 0, 1, 1),
		(drawing, 3469, 3469, 0, 0, 0, 0, 1, 1),
		(drawing, 3468, 3468, 0, 0, 0, 0, 1, 1),
		(drawing, 3467, 3467, 0, 0, 0, 0, 1, 1),
		(drawing, 3466, 3466, 0, 0, 0, 0, 1, 1),
		(drawing, 3465, 3465, 0, 0, 0, 0, 1, 1),
		(drawing, 3464, 3464, 0, 0, 0, 0, 1, 1),
		(drawing, 3463, 3463, 0, 0, 0, 0, 1, 1),
		(drawing, 3462, 3462, 0, 0, 0, 0, 1, 1),
		(drawing, 3461, 3461, 0, 0, 0, 0, 1, 1),
		(drawing, 3460, 3460, 0, 0, 0, 0, 1, 1),
		(drawing, 3459, 3459, 0, 0, 0, 0, 1, 1),
		(drawing, 3458, 3458, 0, 0, 0, 0, 1, 1),
		(drawing, 3457, 3457, 0, 0, 0, 0, 1, 1),
		(drawing, 3456, 3456, 0, 0, 0, 0, 1, 1),
		(drawing, 3455, 3455, 0, 0, 0, 0, 1, 1),
		(drawing, 3454, 3454, 0, 0, 0, 0, 1, 1),
		(drawing, 3453, 3453, 0, 0, 0, 0, 1, 1),
		(drawing, 3452, 3452, 0, 0, 0, 0, 1, 1),
		(drawing, 3451, 3451, 0, 0, 0, 0, 1, 1),
		(drawing, 3450, 3450, 0, 0, 0, 0, 1, 1),
		(drawing, 3449, 3449, 0, 0, 0, 0, 1, 1),
		(drawing, 3448, 3448, 0, 0, 0, 0, 1, 1),
		(drawing, 3447, 3447, 0, 0, 0, 0, 1, 1),
		(drawing, 3446, 3446, 0, 0, 0, 0, 1, 1),
		(drawing, 3445, 3445, 0, 0, 0, 0, 1, 1),
		(drawing, 3444, 3444, 0, 0, 0, 0, 1, 1),
		(drawing, 3443, 3443, 0, 0, 0, 0, 1, 1),
		(drawing, 3442, 3442, 0, 0, 0, 0, 1, 1),
		(drawing, 3441, 3441, 0, 0, 0, 0, 1, 1),
		(drawing, 3440, 3440, 0, 0, 0, 0, 1, 1),
		(drawing, 3439, 3439, 0, 0, 0, 0, 1, 1),
		(drawing, 3438, 3438, 0, 0, 0, 0, 1, 1),
		(drawing, 3437, 3437, 0, 0, 0, 0, 1, 1),
		(drawing, 3436, 3436, 0, 0, 0, 0, 1, 1),
		(drawing, 3435, 3435, 0, 0, 0, 0, 1, 1),
		(drawing, 3434, 3434, 0, 0, 0, 0, 1, 1),
		(drawing, 3433, 3433, 0, 0, 0, 0, 1, 1),
		(drawing, 3432, 3432, 0, 0, 0, 0, 1, 1),
		(drawing, 3431, 3431, 0, 0, 0, 0, 1, 1),
		(drawing, 3430, 3430, 0, 0, 0, 0, 1, 1),
		(drawing, 3429, 3429, 0, 0, 0, 0, 1, 1),
		(drawing, 3428, 3428, 0, 0, 0, 0, 1, 1),
		(drawing, 3427, 3427, 0, 0, 0, 0, 1, 1),
		(drawing, 3426, 3426, 0, 0, 0, 0, 1, 1),
		(drawing, 3425, 3425, 0, 0, 0, 0, 1, 1),
		(drawing, 3424, 3424, 0, 0, 0, 0, 1, 1),
		(drawing, 3423, 3423, 0, 0, 0, 0, 1, 1),
		(drawing, 3422, 3422, 0, 0, 0, 0, 1, 1),
		(drawing, 3421, 3421, 0, 0, 0, 0, 1, 1),
		(drawing, 3420, 3420, 0, 0, 0, 0, 1, 1),
		(drawing, 3419, 3419, 0, 0, 0, 0, 1, 1),
		(drawing, 3418, 3418, 0, 0, 0, 0, 1, 1),
		(drawing, 3417, 3417, 0, 0, 0, 0, 1, 1),
		(drawing, 3416, 3416, 0, 0, 0, 0, 1, 1),
		(drawing, 3415, 3415, 0, 0, 0, 0, 1, 1),
		(drawing, 3414, 3414, 0, 0, 0, 0, 1, 1),
		(drawing, 3413, 3413, 0, 0, 0, 0, 1, 1),
		(drawing, 3412, 3412, 0, 0, 0, 0, 1, 1),
		(drawing, 3411, 3411, 0, 0, 0, 0, 1, 1),
		(drawing, 3410, 3410, 0, 0, 0, 0, 1, 1),
		(drawing, 3409, 3409, 0, 0, 0, 0, 1, 1),
		(drawing, 3408, 3408, 0, 0, 0, 0, 1, 1),
		(drawing, 3407, 3407, 0, 0, 0, 0, 1, 1),
		(drawing, 3406, 3406, 0, 0, 0, 0, 1, 1),
		(drawing, 3405, 3405, 0, 0, 0, 0, 1, 1),
		(drawing, 3404, 3404, 0, 0, 0, 0, 1, 1),
		(drawing, 3403, 3403, 0, 0, 0, 0, 1, 1),
		(drawing, 3402, 3402, 0, 0, 0, 0, 1, 1),
		(drawing, 3401, 3401, 0, 0, 0, 0, 1, 1),
		(drawing, 3400, 3400, 0, 0, 0, 0, 1, 1),
		(drawing, 3399, 3399, 0, 0, 0, 0, 1, 1),
		(drawing, 3398, 3398, 0, 0, 0, 0, 1, 1),
		(drawing, 3397, 3397, 0, 0, 0, 0, 1, 1),
		(drawing, 3396, 3396, 0, 0, 0, 0, 1, 1),
		(drawing, 3395, 3395, 0, 0, 0, 0, 1, 1),
		(drawing, 3394, 3394, 0, 0, 0, 0, 1, 1),
		(drawing, 3393, 3393, 0, 0, 0, 0, 1, 1),
		(drawing, 3392, 3392, 0, 0, 0, 0, 1, 1),
		(drawing, 3391, 3391, 0, 0, 0, 0, 1, 1),
		(drawing, 3390, 3390, 0, 0, 0, 0, 1, 1),
		(drawing, 3389, 3389, 0, 0, 0, 0, 1, 1),
		(drawing, 3388, 3388, 0, 0, 0, 0, 1, 1),
		(drawing, 3387, 3387, 0, 0, 0, 0, 1, 1),
		(drawing, 3386, 3386, 0, 0, 0, 0, 1, 1),
		(drawing, 3385, 3385, 0, 0, 0, 0, 1, 1),
		(drawing, 3384, 3384, 0, 0, 0, 0, 1, 1),
		(drawing, 3383, 3383, 0, 0, 0, 0, 1, 1),
		(drawing, 3382, 3382, 0, 0, 0, 0, 1, 1),
		(drawing, 3381, 3381, 0, 0, 0, 0, 1, 1),
		(drawing, 3380, 3380, 0, 0, 0, 0, 1, 1),
		(drawing, 3379, 3379, 0, 0, 0, 0, 1, 1),
		(drawing, 3378, 3378, 0, 0, 0, 0, 1, 1),
		(drawing, 3377, 3377, 0, 0, 0, 0, 1, 1),
		(drawing, 3376, 3376, 0, 0, 0, 0, 1, 1),
		(drawing, 3375, 3375, 0, 0, 0, 0, 1, 1),
		(drawing, 3374, 3374, 0, 0, 0, 0, 1, 1),
		(drawing, 3373, 3373, 0, 0, 0, 0, 1, 1),
		(drawing, 3372, 3372, 0, 0, 0, 0, 1, 1),
		(drawing, 3371, 3371, 0, 0, 0, 0, 1, 1),
		(drawing, 3370, 3370, 0, 0, 0, 0, 1, 1),
		(drawing, 3369, 3369, 0, 0, 0, 0, 1, 1),
		(drawing, 3368, 3368, 0, 0, 0, 0, 1, 1),
		(drawing, 3367, 3367, 0, 0, 0, 0, 1, 1),
		(drawing, 3366, 3366, 0, 0, 0, 0, 1, 1),
		(drawing, 3365, 3365, 0, 0, 0, 0, 1, 1),
		(drawing, 3364, 3364, 0, 0, 0, 0, 1, 1),
		(drawing, 3363, 3363, 0, 0, 0, 0, 1, 1),
		(drawing, 3362, 3362, 0, 0, 0, 0, 1, 1),
		(drawing, 3361, 3361, 0, 0, 0, 0, 1, 1),
		(drawing, 3360, 3360, 0, 0, 0, 0, 1, 1),
		(drawing, 3359, 3359, 0, 0, 0, 0, 1, 1),
		(drawing, 3358, 3358, 0, 0, 0, 0, 1, 1),
		(drawing, 3357, 3357, 0, 0, 0, 0, 1, 1),
		(drawing, 3356, 3356, 0, 0, 0, 0, 1, 1),
		(drawing, 3355, 3355, 0, 0, 0, 0, 1, 1),
		(drawing, 3354, 3354, 0, 0, 0, 0, 1, 1),
		(drawing, 3353, 3353, 0, 0, 0, 0, 1, 1),
		(drawing, 3352, 3352, 0, 0, 0, 0, 1, 1),
		(drawing, 3351, 3351, 0, 0, 0, 0, 1, 1),
		(drawing, 3350, 3350, 0, 0, 0, 0, 1, 1),
		(drawing, 3349, 3349, 0, 0, 0, 0, 1, 1),
		(drawing, 3348, 3348, 0, 0, 0, 0, 1, 1),
		(drawing, 3347, 3347, 0, 0, 0, 0, 1, 1),
		(drawing, 3346, 3346, 0, 0, 0, 0, 1, 1),
		(drawing, 3345, 3345, 0, 0, 0, 0, 1, 1),
		(drawing, 3344, 3344, 0, 0, 0, 0, 1, 1),
		(drawing, 3343, 3343, 0, 0, 0, 0, 1, 1),
		(drawing, 3342, 3342, 0, 0, 0, 0, 1, 1),
		(drawing, 3341, 3341, 0, 0, 0, 0, 1, 1),
		(drawing, 3340, 3340, 0, 0, 0, 0, 1, 1),
		(drawing, 3339, 3339, 0, 0, 0, 0, 1, 1),
		(drawing, 3338, 3338, 0, 0, 0, 0, 1, 1),
		(drawing, 3337, 3337, 0, 0, 0, 0, 1, 1),
		(drawing, 3336, 3336, 0, 0, 0, 0, 1, 1),
		(drawing, 3335, 3335, 0, 0, 0, 0, 1, 1),
		(drawing, 3334, 3334, 0, 0, 0, 0, 1, 1),
		(drawing, 3333, 3333, 0, 0, 0, 0, 1, 1),
		(drawing, 3332, 3332, 0, 0, 0, 0, 1, 1),
		(drawing, 3331, 3331, 0, 0, 0, 0, 1, 1),
		(drawing, 3330, 3330, 0, 0, 0, 0, 1, 1),
		(drawing, 3329, 3329, 0, 0, 0, 0, 1, 1),
		(drawing, 3328, 3328, 0, 0, 0, 0, 1, 1),
		(drawing, 3327, 3327, 0, 0, 0, 0, 1, 1),
		(drawing, 3326, 3326, 0, 0, 0, 0, 1, 1),
		(drawing, 3325, 3325, 0, 0, 0, 0, 1, 1),
		(drawing, 3324, 3324, 0, 0, 0, 0, 1, 1),
		(drawing, 3323, 3323, 0, 0, 0, 0, 1, 1),
		(drawing, 3322, 3322, 0, 0, 0, 0, 1, 1),
		(drawing, 3321, 3321, 0, 0, 0, 0, 1, 1),
		(drawing, 3320, 3320, 0, 0, 0, 0, 1, 1),
		(drawing, 3319, 3319, 0, 0, 0, 0, 1, 1),
		(drawing, 3318, 3318, 0, 0, 0, 0, 1, 1),
		(drawing, 3317, 3317, 0, 0, 0, 0, 1, 1),
		(drawing, 3316, 3316, 0, 0, 0, 0, 1, 1),
		(drawing, 3315, 3315, 0, 0, 0, 0, 1, 1),
		(drawing, 3314, 3314, 0, 0, 0, 0, 1, 1),
		(drawing, 3313, 3313, 0, 0, 0, 0, 1, 1),
		(drawing, 3312, 3312, 0, 0, 0, 0, 1, 1),
		(drawing, 3311, 3311, 0, 0, 0, 0, 1, 1),
		(drawing, 3310, 3310, 0, 0, 0, 0, 1, 1),
		(drawing, 3309, 3309, 0, 0, 0, 0, 1, 1),
		(drawing, 3308, 3308, 0, 0, 0, 0, 1, 1),
		(drawing, 3307, 3307, 0, 0, 0, 0, 1, 1),
		(drawing, 3306, 3306, 0, 0, 0, 0, 1, 1),
		(drawing, 3305, 3305, 0, 0, 0, 0, 1, 1),
		(drawing, 3304, 3304, 0, 0, 0, 0, 1, 1),
		(drawing, 3303, 3303, 0, 0, 0, 0, 1, 1),
		(drawing, 3302, 3302, 0, 0, 0, 0, 1, 1),
		(drawing, 3301, 3301, 0, 0, 0, 0, 1, 1),
		(drawing, 3300, 3300, 0, 0, 0, 0, 1, 1),
		(drawing, 3299, 3299, 0, 0, 0, 0, 1, 1),
		(drawing, 3298, 3298, 0, 0, 0, 0, 1, 1),
		(drawing, 3297, 3297, 0, 0, 0, 0, 1, 1),
		(drawing, 3296, 3296, 0, 0, 0, 0, 1, 1),
		(drawing, 3295, 3295, 0, 0, 0, 0, 1, 1),
		(drawing, 3294, 3294, 0, 0, 0, 0, 1, 1),
		(drawing, 3293, 3293, 0, 0, 0, 0, 1, 1),
		(drawing, 3292, 3292, 0, 0, 0, 0, 1, 1),
		(drawing, 3291, 3291, 0, 0, 0, 0, 1, 1),
		(drawing, 3290, 3290, 0, 0, 0, 0, 1, 1),
		(drawing, 3289, 3289, 0, 0, 0, 0, 1, 1),
		(drawing, 3288, 3288, 0, 0, 0, 0, 1, 1),
		(drawing, 3287, 3287, 0, 0, 0, 0, 1, 1),
		(drawing, 3286, 3286, 0, 0, 0, 0, 1, 1),
		(drawing, 3285, 3285, 0, 0, 0, 0, 1, 1),
		(drawing, 3284, 3284, 0, 0, 0, 0, 1, 1),
		(drawing, 3283, 3283, 0, 0, 0, 0, 1, 1),
		(drawing, 3282, 3282, 0, 0, 0, 0, 1, 1),
		(drawing, 3281, 3281, 0, 0, 0, 0, 1, 1),
		(drawing, 3280, 3280, 0, 0, 0, 0, 1, 1),
		(drawing, 3279, 3279, 0, 0, 0, 0, 1, 1),
		(drawing, 3278, 3278, 0, 0, 0, 0, 1, 1),
		(drawing, 3277, 3277, 0, 0, 0, 0, 1, 1),
		(drawing, 3276, 3276, 0, 0, 0, 0, 1, 1),
		(drawing, 3275, 3275, 0, 0, 0, 0, 1, 1),
		(drawing, 3274, 3274, 0, 0, 0, 0, 1, 1),
		(drawing, 3273, 3273, 0, 0, 0, 0, 1, 1),
		(drawing, 3272, 3272, 0, 0, 0, 0, 1, 1),
		(drawing, 3271, 3271, 0, 0, 0, 0, 1, 1),
		(drawing, 3270, 3270, 0, 0, 0, 0, 1, 1),
		(drawing, 3269, 3269, 0, 0, 0, 0, 1, 1),
		(drawing, 3268, 3268, 0, 0, 0, 0, 1, 1),
		(drawing, 3267, 3267, 0, 0, 0, 0, 1, 1),
		(drawing, 3266, 3266, 0, 0, 0, 0, 1, 1),
		(drawing, 3265, 3265, 0, 0, 0, 0, 1, 1),
		(drawing, 3264, 3264, 0, 0, 0, 0, 1, 1),
		(drawing, 3263, 3263, 0, 0, 0, 0, 1, 1),
		(drawing, 3262, 3262, 0, 0, 0, 0, 1, 1),
		(drawing, 3261, 3261, 0, 0, 0, 0, 1, 1),
		(drawing, 3260, 3260, 0, 0, 0, 0, 1, 1),
		(drawing, 3259, 3259, 0, 0, 0, 0, 1, 1),
		(drawing, 3258, 3258, 0, 0, 0, 0, 1, 1),
		(drawing, 3257, 3257, 0, 0, 0, 0, 1, 1),
		(drawing, 3256, 3256, 0, 0, 0, 0, 1, 1),
		(drawing, 3255, 3255, 0, 0, 0, 0, 1, 1),
		(drawing, 3254, 3254, 0, 0, 0, 0, 1, 1),
		(drawing, 3253, 3253, 0, 0, 0, 0, 1, 1),
		(drawing, 3252, 3252, 0, 0, 0, 0, 1, 1),
		(drawing, 3251, 3251, 0, 0, 0, 0, 1, 1),
		(drawing, 3250, 3250, 0, 0, 0, 0, 1, 1),
		(drawing, 3249, 3249, 0, 0, 0, 0, 1, 1),
		(drawing, 3248, 3248, 0, 0, 0, 0, 1, 1),
		(drawing, 3247, 3247, 0, 0, 0, 0, 1, 1),
		(drawing, 3246, 3246, 0, 0, 0, 0, 1, 1),
		(drawing, 3245, 3245, 0, 0, 0, 0, 1, 1),
		(drawing, 3244, 3244, 0, 0, 0, 0, 1, 1),
		(drawing, 3243, 3243, 0, 0, 0, 0, 1, 1),
		(drawing, 3242, 3242, 0, 0, 0, 0, 1, 1),
		(drawing, 3241, 3241, 0, 0, 0, 0, 1, 1),
		(drawing, 3240, 3240, 0, 0, 0, 0, 1, 1),
		(drawing, 3239, 3239, 0, 0, 0, 0, 1, 1),
		(drawing, 3238, 3238, 0, 0, 0, 0, 1, 1),
		(drawing, 3237, 3237, 0, 0, 0, 0, 1, 1),
		(drawing, 3236, 3236, 0, 0, 0, 0, 1, 1),
		(drawing, 3235, 3235, 0, 0, 0, 0, 1, 1),
		(drawing, 3234, 3234, 0, 0, 0, 0, 1, 1),
		(drawing, 3233, 3233, 0, 0, 0, 0, 1, 1),
		(drawing, 3232, 3232, 0, 0, 0, 0, 1, 1),
		(drawing, 3231, 3231, 0, 0, 0, 0, 1, 1),
		(drawing, 3230, 3230, 0, 0, 0, 0, 1, 1),
		(drawing, 3229, 3229, 0, 0, 0, 0, 1, 1),
		(drawing, 3228, 3228, 0, 0, 0, 0, 1, 1),
		(drawing, 3227, 3227, 0, 0, 0, 0, 1, 1),
		(drawing, 3226, 3226, 0, 0, 0, 0, 1, 1),
		(drawing, 3225, 3225, 0, 0, 0, 0, 1, 1),
		(drawing, 3224, 3224, 0, 0, 0, 0, 1, 1),
		(drawing, 3223, 3223, 0, 0, 0, 0, 1, 1),
		(drawing, 3222, 3222, 0, 0, 0, 0, 1, 1),
		(drawing, 3221, 3221, 0, 0, 0, 0, 1, 1),
		(drawing, 3220, 3220, 0, 0, 0, 0, 1, 1),
		(drawing, 3219, 3219, 0, 0, 0, 0, 1, 1),
		(drawing, 3218, 3218, 0, 0, 0, 0, 1, 1),
		(drawing, 3217, 3217, 0, 0, 0, 0, 1, 1),
		(drawing, 3216, 3216, 0, 0, 0, 0, 1, 1),
		(drawing, 3215, 3215, 0, 0, 0, 0, 1, 1),
		(drawing, 3214, 3214, 0, 0, 0, 0, 1, 1),
		(drawing, 3213, 3213, 0, 0, 0, 0, 1, 1),
		(drawing, 3212, 3212, 0, 0, 0, 0, 1, 1),
		(drawing, 3211, 3211, 0, 0, 0, 0, 1, 1),
		(drawing, 3210, 3210, 0, 0, 0, 0, 1, 1),
		(drawing, 3209, 3209, 0, 0, 0, 0, 1, 1),
		(drawing, 3208, 3208, 0, 0, 0, 0, 1, 1),
		(drawing, 3207, 3207, 0, 0, 0, 0, 1, 1),
		(drawing, 3206, 3206, 0, 0, 0, 0, 1, 1),
		(drawing, 3205, 3205, 0, 0, 0, 0, 1, 1),
		(drawing, 3204, 3204, 0, 0, 0, 0, 1, 1),
		(drawing, 3203, 3203, 0, 0, 0, 0, 1, 1),
		(drawing, 3202, 3202, 0, 0, 0, 0, 1, 1),
		(drawing, 3201, 3201, 0, 0, 0, 0, 1, 1),
		(drawing, 3200, 3200, 0, 0, 0, 0, 1, 1),
		(drawing, 3199, 3199, 0, 0, 0, 0, 1, 1),
		(drawing, 3198, 3198, 0, 0, 0, 0, 1, 1),
		(drawing, 3197, 3197, 0, 0, 0, 0, 1, 1),
		(drawing, 3196, 3196, 0, 0, 0, 0, 1, 1),
		(drawing, 3195, 3195, 0, 0, 0, 0, 1, 1),
		(drawing, 3194, 3194, 0, 0, 0, 0, 1, 1),
		(drawing, 3193, 3193, 0, 0, 0, 0, 1, 1),
		(drawing, 3192, 3192, 0, 0, 0, 0, 1, 1),
		(drawing, 3191, 3191, 0, 0, 0, 0, 1, 1),
		(drawing, 3190, 3190, 0, 0, 0, 0, 1, 1),
		(drawing, 3189, 3189, 0, 0, 0, 0, 1, 1),
		(drawing, 3188, 3188, 0, 0, 0, 0, 1, 1),
		(drawing, 3187, 3187, 0, 0, 0, 0, 1, 1),
		(drawing, 3186, 3186, 0, 0, 0, 0, 1, 1),
		(drawing, 3185, 3185, 0, 0, 0, 0, 1, 1),
		(drawing, 3184, 3184, 0, 0, 0, 0, 1, 1),
		(drawing, 3183, 3183, 0, 0, 0, 0, 1, 1),
		(drawing, 3182, 3182, 0, 0, 0, 0, 1, 1),
		(drawing, 3181, 3181, 0, 0, 0, 0, 1, 1),
		(drawing, 3180, 3180, 0, 0, 0, 0, 1, 1),
		(drawing, 3179, 3179, 0, 0, 0, 0, 1, 1),
		(drawing, 3178, 3178, 0, 0, 0, 0, 1, 1),
		(drawing, 3177, 3177, 0, 0, 0, 0, 1, 1),
		(drawing, 3176, 3176, 0, 0, 0, 0, 1, 1),
		(drawing, 3175, 3175, 0, 0, 0, 0, 1, 1),
		(drawing, 3174, 3174, 0, 0, 0, 0, 1, 1),
		(drawing, 3173, 3173, 0, 0, 0, 0, 1, 1),
		(drawing, 3172, 3172, 0, 0, 0, 0, 1, 1),
		(drawing, 3171, 3171, 0, 0, 0, 0, 1, 1),
		(drawing, 3170, 3170, 0, 0, 0, 0, 1, 1),
		(drawing, 3169, 3169, 0, 0, 0, 0, 1, 1),
		(drawing, 3168, 3168, 0, 0, 0, 0, 1, 1),
		(drawing, 3167, 3167, 0, 0, 0, 0, 1, 1),
		(drawing, 3166, 3166, 0, 0, 0, 0, 1, 1),
		(drawing, 3165, 3165, 0, 0, 0, 0, 1, 1),
		(drawing, 3164, 3164, 0, 0, 0, 0, 1, 1),
		(drawing, 3163, 3163, 0, 0, 0, 0, 1, 1),
		(drawing, 3162, 3162, 0, 0, 0, 0, 1, 1),
		(drawing, 3161, 3161, 0, 0, 0, 0, 1, 1),
		(drawing, 3160, 3160, 0, 0, 0, 0, 1, 1),
		(drawing, 3159, 3159, 0, 0, 0, 0, 1, 1),
		(drawing, 3158, 3158, 0, 0, 0, 0, 1, 1),
		(drawing, 3157, 3157, 0, 0, 0, 0, 1, 1),
		(drawing, 3156, 3156, 0, 0, 0, 0, 1, 1),
		(drawing, 3155, 3155, 0, 0, 0, 0, 1, 1),
		(drawing, 3154, 3154, 0, 0, 0, 0, 1, 1),
		(drawing, 3153, 3153, 0, 0, 0, 0, 1, 1),
		(drawing, 3152, 3152, 0, 0, 0, 0, 1, 1),
		(drawing, 3151, 3151, 0, 0, 0, 0, 1, 1),
		(drawing, 3150, 3150, 0, 0, 0, 0, 1, 1),
		(drawing, 3149, 3149, 0, 0, 0, 0, 1, 1),
		(drawing, 3148, 3148, 0, 0, 0, 0, 1, 1),
		(drawing, 3147, 3147, 0, 0, 0, 0, 1, 1),
		(drawing, 3146, 3146, 0, 0, 0, 0, 1, 1),
		(drawing, 3145, 3145, 0, 0, 0, 0, 1, 1),
		(drawing, 3144, 3144, 0, 0, 0, 0, 1, 1),
		(drawing, 3143, 3143, 0, 0, 0, 0, 1, 1),
		(drawing, 3142, 3142, 0, 0, 0, 0, 1, 1),
		(drawing, 3141, 3141, 0, 0, 0, 0, 1, 1),
		(drawing, 3140, 3140, 0, 0, 0, 0, 1, 1),
		(drawing, 3139, 3139, 0, 0, 0, 0, 1, 1),
		(drawing, 3138, 3138, 0, 0, 0, 0, 1, 1),
		(drawing, 3137, 3137, 0, 0, 0, 0, 1, 1),
		(drawing, 3136, 3136, 0, 0, 0, 0, 1, 1),
		(drawing, 3135, 3135, 0, 0, 0, 0, 1, 1),
		(drawing, 3134, 3134, 0, 0, 0, 0, 1, 1),
		(drawing, 3133, 3133, 0, 0, 0, 0, 1, 1),
		(drawing, 3132, 3132, 0, 0, 0, 0, 1, 1),
		(drawing, 3131, 3131, 0, 0, 0, 0, 1, 1),
		(drawing, 3130, 3130, 0, 0, 0, 0, 1, 1),
		(drawing, 3129, 3129, 0, 0, 0, 0, 1, 1),
		(drawing, 3128, 3128, 0, 0, 0, 0, 1, 1),
		(drawing, 3127, 3127, 0, 0, 0, 0, 1, 1),
		(drawing, 3126, 3126, 0, 0, 0, 0, 1, 1),
		(drawing, 3125, 3125, 0, 0, 0, 0, 1, 1),
		(drawing, 3124, 3124, 0, 0, 0, 0, 1, 1),
		(drawing, 3123, 3123, 0, 0, 0, 0, 1, 1),
		(drawing, 3122, 3122, 0, 0, 0, 0, 1, 1),
		(drawing, 3121, 3121, 0, 0, 0, 0, 1, 1),
		(drawing, 3120, 3120, 0, 0, 0, 0, 1, 1),
		(drawing, 3119, 3119, 0, 0, 0, 0, 1, 1),
		(drawing, 3118, 3118, 0, 0, 0, 0, 1, 1),
		(drawing, 3117, 3117, 0, 0, 0, 0, 1, 1),
		(drawing, 3116, 3116, 0, 0, 0, 0, 1, 1),
		(drawing, 3115, 3115, 0, 0, 0, 0, 1, 1),
		(drawing, 3114, 3114, 0, 0, 0, 0, 1, 1),
		(drawing, 3113, 3113, 0, 0, 0, 0, 1, 1),
		(drawing, 3112, 3112, 0, 0, 0, 0, 1, 1),
		(drawing, 3111, 3111, 0, 0, 0, 0, 1, 1),
		(drawing, 3110, 3110, 0, 0, 0, 0, 1, 1),
		(drawing, 3109, 3109, 0, 0, 0, 0, 1, 1),
		(drawing, 3108, 3108, 0, 0, 0, 0, 1, 1),
		(drawing, 3107, 3107, 0, 0, 0, 0, 1, 1),
		(drawing, 3106, 3106, 0, 0, 0, 0, 1, 1),
		(drawing, 3105, 3105, 0, 0, 0, 0, 1, 1),
		(drawing, 3104, 3104, 0, 0, 0, 0, 1, 1),
		(drawing, 3103, 3103, 0, 0, 0, 0, 1, 1),
		(drawing, 3102, 3102, 0, 0, 0, 0, 1, 1),
		(drawing, 3101, 3101, 0, 0, 0, 0, 1, 1),
		(drawing, 3100, 3100, 0, 0, 0, 0, 1, 1),
		(drawing, 3099, 3099, 0, 0, 0, 0, 1, 1),
		(drawing, 3098, 3098, 0, 0, 0, 0, 1, 1),
		(drawing, 3097, 3097, 0, 0, 0, 0, 1, 1),
		(drawing, 3096, 3096, 0, 0, 0, 0, 1, 1),
		(drawing, 3095, 3095, 0, 0, 0, 0, 1, 1),
		(drawing, 3094, 3094, 0, 0, 0, 0, 1, 1),
		(drawing, 3093, 3093, 0, 0, 0, 0, 1, 1),
		(drawing, 3092, 3092, 0, 0, 0, 0, 1, 1),
		(drawing, 3091, 3091, 0, 0, 0, 0, 1, 1),
		(drawing, 3090, 3090, 0, 0, 0, 0, 1, 1),
		(drawing, 3089, 3089, 0, 0, 0, 0, 1, 1),
		(drawing, 3088, 3088, 0, 0, 0, 0, 1, 1),
		(drawing, 3087, 3087, 0, 0, 0, 0, 1, 1),
		(drawing, 3086, 3086, 0, 0, 0, 0, 1, 1),
		(drawing, 3085, 3085, 0, 0, 0, 0, 1, 1),
		(drawing, 3084, 3084, 0, 0, 0, 0, 1, 1),
		(drawing, 3083, 3083, 0, 0, 0, 0, 1, 1),
		(drawing, 3082, 3082, 0, 0, 0, 0, 1, 1),
		(drawing, 3081, 3081, 0, 0, 0, 0, 1, 1),
		(drawing, 3080, 3080, 0, 0, 0, 0, 1, 1),
		(drawing, 3079, 3079, 0, 0, 0, 0, 1, 1),
		(drawing, 3078, 3078, 0, 0, 0, 0, 1, 1),
		(drawing, 3077, 3077, 0, 0, 0, 0, 1, 1),
		(drawing, 3076, 3076, 0, 0, 0, 0, 1, 1),
		(drawing, 3075, 3075, 0, 0, 0, 0, 1, 1),
		(drawing, 3074, 3074, 0, 0, 0, 0, 1, 1),
		(drawing, 3073, 3073, 0, 0, 0, 0, 1, 1),
		(drawing, 3072, 3072, 0, 0, 0, 0, 1, 1),
		(drawing, 3071, 3071, 0, 0, 0, 0, 1, 1),
		(drawing, 3070, 3070, 0, 0, 0, 0, 1, 1),
		(drawing, 3069, 3069, 0, 0, 0, 0, 1, 1),
		(drawing, 3068, 3068, 0, 0, 0, 0, 1, 1),
		(drawing, 3067, 3067, 0, 0, 0, 0, 1, 1),
		(drawing, 3066, 3066, 0, 0, 0, 0, 1, 1),
		(drawing, 3065, 3065, 0, 0, 0, 0, 1, 1),
		(drawing, 3064, 3064, 0, 0, 0, 0, 1, 1),
		(drawing, 3063, 3063, 0, 0, 0, 0, 1, 1),
		(drawing, 3062, 3062, 0, 0, 0, 0, 1, 1),
		(drawing, 3061, 3061, 0, 0, 0, 0, 1, 1),
		(drawing, 3060, 3060, 0, 0, 0, 0, 1, 1),
		(drawing, 3059, 3059, 0, 0, 0, 0, 1, 1),
		(drawing, 3058, 3058, 0, 0, 0, 0, 1, 1),
		(drawing, 3057, 3057, 0, 0, 0, 0, 1, 1),
		(drawing, 3056, 3056, 0, 0, 0, 0, 1, 1),
		(drawing, 3055, 3055, 0, 0, 0, 0, 1, 1),
		(drawing, 3054, 3054, 0, 0, 0, 0, 1, 1),
		(drawing, 3053, 3053, 0, 0, 0, 0, 1, 1),
		(drawing, 3052, 3052, 0, 0, 0, 0, 1, 1),
		(drawing, 3051, 3051, 0, 0, 0, 0, 1, 1),
		(drawing, 3050, 3050, 0, 0, 0, 0, 1, 1),
		(drawing, 3049, 3049, 0, 0, 0, 0, 1, 1),
		(drawing, 3048, 3048, 0, 0, 0, 0, 1, 1),
		(drawing, 3047, 3047, 0, 0, 0, 0, 1, 1),
		(drawing, 3046, 3046, 0, 0, 0, 0, 1, 1),
		(drawing, 3045, 3045, 0, 0, 0, 0, 1, 1),
		(drawing, 3044, 3044, 0, 0, 0, 0, 1, 1),
		(drawing, 3043, 3043, 0, 0, 0, 0, 1, 1),
		(drawing, 3042, 3042, 0, 0, 0, 0, 1, 1),
		(drawing, 3041, 3041, 0, 0, 0, 0, 1, 1),
		(drawing, 3040, 3040, 0, 0, 0, 0, 1, 1),
		(drawing, 3039, 3039, 0, 0, 0, 0, 1, 1),
		(drawing, 3038, 3038, 0, 0, 0, 0, 1, 1),
		(drawing, 3037, 3037, 0, 0, 0, 0, 1, 1),
		(drawing, 3036, 3036, 0, 0, 0, 0, 1, 1),
		(drawing, 3035, 3035, 0, 0, 0, 0, 1, 1),
		(drawing, 3034, 3034, 0, 0, 0, 0, 1, 1),
		(drawing, 3033, 3033, 0, 0, 0, 0, 1, 1),
		(drawing, 3032, 3032, 0, 0, 0, 0, 1, 1),
		(drawing, 3031, 3031, 0, 0, 0, 0, 1, 1),
		(drawing, 3030, 3030, 0, 0, 0, 0, 1, 1),
		(drawing, 3029, 3029, 0, 0, 0, 0, 1, 1),
		(drawing, 3028, 3028, 0, 0, 0, 0, 1, 1),
		(drawing, 3027, 3027, 0, 0, 0, 0, 1, 1),
		(drawing, 3026, 3026, 0, 0, 0, 0, 1, 1),
		(drawing, 3025, 3025, 0, 0, 0, 0, 1, 1),
		(drawing, 3024, 3024, 0, 0, 0, 0, 1, 1),
		(drawing, 3023, 3023, 0, 0, 0, 0, 1, 1),
		(drawing, 3022, 3022, 0, 0, 0, 0, 1, 1),
		(drawing, 3021, 3021, 0, 0, 0, 0, 1, 1),
		(drawing, 3020, 3020, 0, 0, 0, 0, 1, 1),
		(drawing, 3019, 3019, 0, 0, 0, 0, 1, 1),
		(drawing, 3018, 3018, 0, 0, 0, 0, 1, 1),
		(drawing, 3017, 3017, 0, 0, 0, 0, 1, 1),
		(drawing, 3016, 3016, 0, 0, 0, 0, 1, 1),
		(drawing, 3015, 3015, 0, 0, 0, 0, 1, 1),
		(drawing, 3014, 3014, 0, 0, 0, 0, 1, 1),
		(drawing, 3013, 3013, 0, 0, 0, 0, 1, 1),
		(drawing, 3012, 3012, 0, 0, 0, 0, 1, 1),
		(drawing, 3011, 3011, 0, 0, 0, 0, 1, 1),
		(drawing, 3010, 3010, 0, 0, 0, 0, 1, 1),
		(drawing, 3009, 3009, 0, 0, 0, 0, 1, 1),
		(drawing, 3008, 3008, 0, 0, 0, 0, 1, 1),
		(drawing, 3007, 3007, 0, 0, 0, 0, 1, 1),
		(drawing, 3006, 3006, 0, 0, 0, 0, 1, 1),
		(drawing, 3005, 3005, 0, 0, 0, 0, 1, 1),
		(drawing, 3004, 3004, 0, 0, 0, 0, 1, 1),
		(drawing, 3003, 3003, 0, 0, 0, 0, 1, 1),
		(drawing, 3002, 3002, 0, 0, 0, 0, 1, 1),
		(drawing, 3001, 3001, 0, 0, 0, 0, 1, 1),
		(drawing, 3000, 3000, 0, 0, 0, 0, 1, 1),
		(drawing, 2999, 2999, 0, 0, 0, 0, 1, 1),
		(drawing, 2998, 2998, 0, 0, 0, 0, 1, 1),
		(drawing, 2997, 2997, 0, 0, 0, 0, 1, 1),
		(drawing, 2996, 2996, 0, 0, 0, 0, 1, 1),
		(drawing, 2995, 2995, 0, 0, 0, 0, 1, 1),
		(drawing, 2994, 2994, 0, 0, 0, 0, 1, 1),
		(drawing, 2993, 2993, 0, 0, 0, 0, 1, 1),
		(drawing, 2992, 2992, 0, 0, 0, 0, 1, 1),
		(drawing, 2991, 2991, 0, 0, 0, 0, 1, 1),
		(drawing, 2990, 2990, 0, 0, 0, 0, 1, 1),
		(drawing, 2989, 2989, 0, 0, 0, 0, 1, 1),
		(drawing, 2988, 2988, 0, 0, 0, 0, 1, 1),
		(drawing, 2987, 2987, 0, 0, 0, 0, 1, 1),
		(drawing, 2986, 2986, 0, 0, 0, 0, 1, 1),
		(drawing, 2985, 2985, 0, 0, 0, 0, 1, 1),
		(drawing, 2984, 2984, 0, 0, 0, 0, 1, 1),
		(drawing, 2983, 2983, 0, 0, 0, 0, 1, 1),
		(drawing, 2982, 2982, 0, 0, 0, 0, 1, 1),
		(drawing, 2981, 2981, 0, 0, 0, 0, 1, 1),
		(drawing, 2980, 2980, 0, 0, 0, 0, 1, 1),
		(drawing, 2979, 2979, 0, 0, 0, 0, 1, 1),
		(drawing, 2978, 2978, 0, 0, 0, 0, 1, 1),
		(drawing, 2977, 2977, 0, 0, 0, 0, 1, 1),
		(drawing, 2976, 2976, 0, 0, 0, 0, 1, 1),
		(drawing, 2975, 2975, 0, 0, 0, 0, 1, 1),
		(drawing, 2974, 2974, 0, 0, 0, 0, 1, 1),
		(drawing, 2973, 2973, 0, 0, 0, 0, 1, 1),
		(drawing, 2972, 2972, 0, 0, 0, 0, 1, 1),
		(drawing, 2971, 2971, 0, 0, 0, 0, 1, 1),
		(drawing, 2970, 2970, 0, 0, 0, 0, 1, 1),
		(drawing, 2969, 2969, 0, 0, 0, 0, 1, 1),
		(drawing, 2968, 2968, 0, 0, 0, 0, 1, 1),
		(drawing, 2967, 2967, 0, 0, 0, 0, 1, 1),
		(drawing, 2966, 2966, 0, 0, 0, 0, 1, 1),
		(drawing, 2965, 2965, 0, 0, 0, 0, 1, 1),
		(drawing, 2964, 2964, 0, 0, 0, 0, 1, 1),
		(drawing, 2963, 2963, 0, 0, 0, 0, 1, 1),
		(drawing, 2962, 2962, 0, 0, 0, 0, 1, 1),
		(drawing, 2961, 2961, 0, 0, 0, 0, 1, 1),
		(drawing, 2960, 2960, 0, 0, 0, 0, 1, 1),
		(drawing, 2959, 2959, 0, 0, 0, 0, 1, 1),
		(drawing, 2958, 2958, 0, 0, 0, 0, 1, 1),
		(drawing, 2957, 2957, 0, 0, 0, 0, 1, 1),
		(drawing, 2956, 2956, 0, 0, 0, 0, 1, 1),
		(drawing, 2955, 2955, 0, 0, 0, 0, 1, 1),
		(drawing, 2954, 2954, 0, 0, 0, 0, 1, 1),
		(drawing, 2953, 2953, 0, 0, 0, 0, 1, 1),
		(drawing, 2952, 2952, 0, 0, 0, 0, 1, 1),
		(drawing, 2951, 2951, 0, 0, 0, 0, 1, 1),
		(drawing, 2950, 2950, 0, 0, 0, 0, 1, 1),
		(drawing, 2949, 2949, 0, 0, 0, 0, 1, 1),
		(drawing, 2948, 2948, 0, 0, 0, 0, 1, 1),
		(drawing, 2947, 2947, 0, 0, 0, 0, 1, 1),
		(drawing, 2946, 2946, 0, 0, 0, 0, 1, 1),
		(drawing, 2945, 2945, 0, 0, 0, 0, 1, 1),
		(drawing, 2944, 2944, 0, 0, 0, 0, 1, 1),
		(drawing, 2943, 2943, 0, 0, 0, 0, 1, 1),
		(drawing, 2942, 2942, 0, 0, 0, 0, 1, 1),
		(drawing, 2941, 2941, 0, 0, 0, 0, 1, 1),
		(drawing, 2940, 2940, 0, 0, 0, 0, 1, 1),
		(drawing, 2939, 2939, 0, 0, 0, 0, 1, 1),
		(drawing, 2938, 2938, 0, 0, 0, 0, 1, 1),
		(drawing, 2937, 2937, 0, 0, 0, 0, 1, 1),
		(drawing, 2936, 2936, 0, 0, 0, 0, 1, 1),
		(drawing, 2935, 2935, 0, 0, 0, 0, 1, 1),
		(drawing, 2934, 2934, 0, 0, 0, 0, 1, 1),
		(drawing, 2933, 2933, 0, 0, 0, 0, 1, 1),
		(drawing, 2932, 2932, 0, 0, 0, 0, 1, 1),
		(drawing, 2931, 2931, 0, 0, 0, 0, 1, 1),
		(drawing, 2930, 2930, 0, 0, 0, 0, 1, 1),
		(drawing, 2929, 2929, 0, 0, 0, 0, 1, 1),
		(drawing, 2928, 2928, 0, 0, 0, 0, 1, 1),
		(drawing, 2927, 2927, 0, 0, 0, 0, 1, 1),
		(drawing, 2926, 2926, 0, 0, 0, 0, 1, 1),
		(drawing, 2925, 2925, 0, 0, 0, 0, 1, 1),
		(drawing, 2924, 2924, 0, 0, 0, 0, 1, 1),
		(drawing, 2923, 2923, 0, 0, 0, 0, 1, 1),
		(drawing, 2922, 2922, 0, 0, 0, 0, 1, 1),
		(drawing, 2921, 2921, 0, 0, 0, 0, 1, 1),
		(drawing, 2920, 2920, 0, 0, 0, 0, 1, 1),
		(drawing, 2919, 2919, 0, 0, 0, 0, 1, 1),
		(drawing, 2918, 2918, 0, 0, 0, 0, 1, 1),
		(drawing, 2917, 2917, 0, 0, 0, 0, 1, 1),
		(drawing, 2916, 2916, 0, 0, 0, 0, 1, 1),
		(drawing, 2915, 2915, 0, 0, 0, 0, 1, 1),
		(drawing, 2914, 2914, 0, 0, 0, 0, 1, 1),
		(drawing, 2913, 2913, 0, 0, 0, 0, 1, 1),
		(drawing, 2912, 2912, 0, 0, 0, 0, 1, 1),
		(drawing, 2911, 2911, 0, 0, 0, 0, 1, 1),
		(drawing, 2910, 2910, 0, 0, 0, 0, 1, 1),
		(drawing, 2909, 2909, 0, 0, 0, 0, 1, 1),
		(drawing, 2908, 2908, 0, 0, 0, 0, 1, 1),
		(drawing, 2907, 2907, 0, 0, 0, 0, 1, 1),
		(drawing, 2906, 2906, 0, 0, 0, 0, 1, 1),
		(drawing, 2905, 2905, 0, 0, 0, 0, 1, 1),
		(drawing, 2904, 2904, 0, 0, 0, 0, 1, 1),
		(drawing, 2903, 2903, 0, 0, 0, 0, 1, 1),
		(drawing, 2902, 2902, 0, 0, 0, 0, 1, 1),
		(drawing, 2901, 2901, 0, 0, 0, 0, 1, 1),
		(drawing, 2900, 2900, 0, 0, 0, 0, 1, 1),
		(drawing, 2899, 2899, 0, 0, 0, 0, 1, 1),
		(drawing, 2898, 2898, 0, 0, 0, 0, 1, 1),
		(drawing, 2897, 2897, 0, 0, 0, 0, 1, 1),
		(drawing, 2896, 2896, 0, 0, 0, 0, 1, 1),
		(drawing, 2895, 2895, 0, 0, 0, 0, 1, 1),
		(drawing, 2894, 2894, 0, 0, 0, 0, 1, 1),
		(drawing, 2893, 2893, 0, 0, 0, 0, 1, 1),
		(drawing, 2892, 2892, 0, 0, 0, 0, 1, 1),
		(drawing, 2891, 2891, 0, 0, 0, 0, 1, 1),
		(drawing, 2890, 2890, 0, 0, 0, 0, 1, 1),
		(drawing, 2889, 2889, 0, 0, 0, 0, 1, 1),
		(drawing, 2888, 2888, 0, 0, 0, 0, 1, 1),
		(drawing, 2887, 2887, 0, 0, 0, 0, 1, 1),
		(drawing, 2886, 2886, 0, 0, 0, 0, 1, 1),
		(drawing, 2885, 2885, 0, 0, 0, 0, 1, 1),
		(drawing, 2884, 2884, 0, 0, 0, 0, 1, 1),
		(drawing, 2883, 2883, 0, 0, 0, 0, 1, 1),
		(drawing, 2882, 2882, 0, 0, 0, 0, 1, 1),
		(drawing, 2881, 2881, 0, 0, 0, 0, 1, 1),
		(drawing, 2880, 2880, 0, 0, 0, 0, 1, 1),
		(drawing, 2879, 2879, 0, 0, 0, 0, 1, 1),
		(drawing, 2878, 2878, 0, 0, 0, 0, 1, 1),
		(drawing, 2877, 2877, 0, 0, 0, 0, 1, 1),
		(drawing, 2876, 2876, 0, 0, 0, 0, 1, 1),
		(drawing, 2875, 2875, 0, 0, 0, 0, 1, 1),
		(drawing, 2874, 2874, 0, 0, 0, 0, 1, 1),
		(drawing, 2873, 2873, 0, 0, 0, 0, 1, 1),
		(drawing, 2872, 2872, 0, 0, 0, 0, 1, 1),
		(drawing, 2871, 2871, 0, 0, 0, 0, 1, 1),
		(drawing, 2870, 2870, 0, 0, 0, 0, 1, 1),
		(drawing, 2869, 2869, 0, 0, 0, 0, 1, 1),
		(drawing, 2868, 2868, 0, 0, 0, 0, 1, 1),
		(drawing, 2867, 2867, 0, 0, 0, 0, 1, 1),
		(drawing, 2866, 2866, 0, 0, 0, 0, 1, 1),
		(drawing, 2865, 2865, 0, 0, 0, 0, 1, 1),
		(drawing, 2864, 2864, 0, 0, 0, 0, 1, 1),
		(drawing, 2863, 2863, 0, 0, 0, 0, 1, 1),
		(drawing, 2862, 2862, 0, 0, 0, 0, 1, 1),
		(drawing, 2861, 2861, 0, 0, 0, 0, 1, 1),
		(drawing, 2860, 2860, 0, 0, 0, 0, 1, 1),
		(drawing, 2859, 2859, 0, 0, 0, 0, 1, 1),
		(drawing, 2858, 2858, 0, 0, 0, 0, 1, 1),
		(drawing, 2857, 2857, 0, 0, 0, 0, 1, 1),
		(drawing, 2856, 2856, 0, 0, 0, 0, 1, 1),
		(drawing, 2855, 2855, 0, 0, 0, 0, 1, 1),
		(drawing, 2854, 2854, 0, 0, 0, 0, 1, 1),
		(drawing, 2853, 2853, 0, 0, 0, 0, 1, 1),
		(drawing, 2852, 2852, 0, 0, 0, 0, 1, 1),
		(drawing, 2851, 2851, 0, 0, 0, 0, 1, 1),
		(drawing, 2850, 2850, 0, 0, 0, 0, 1, 1),
		(drawing, 2849, 2849, 0, 0, 0, 0, 1, 1),
		(drawing, 2848, 2848, 0, 0, 0, 0, 1, 1),
		(drawing, 2847, 2847, 0, 0, 0, 0, 1, 1),
		(drawing, 2846, 2846, 0, 0, 0, 0, 1, 1),
		(drawing, 2845, 2845, 0, 0, 0, 0, 1, 1),
		(drawing, 2844, 2844, 0, 0, 0, 0, 1, 1),
		(drawing, 2843, 2843, 0, 0, 0, 0, 1, 1),
		(drawing, 2842, 2842, 0, 0, 0, 0, 1, 1),
		(drawing, 2841, 2841, 0, 0, 0, 0, 1, 1),
		(drawing, 2840, 2840, 0, 0, 0, 0, 1, 1),
		(drawing, 2839, 2839, 0, 0, 0, 0, 1, 1),
		(drawing, 2838, 2838, 0, 0, 0, 0, 1, 1),
		(drawing, 2837, 2837, 0, 0, 0, 0, 1, 1),
		(drawing, 2836, 2836, 0, 0, 0, 0, 1, 1),
		(drawing, 2835, 2835, 0, 0, 0, 0, 1, 1),
		(drawing, 2834, 2834, 0, 0, 0, 0, 1, 1),
		(drawing, 2833, 2833, 0, 0, 0, 0, 1, 1),
		(drawing, 2832, 2832, 0, 0, 0, 0, 1, 1),
		(drawing, 2831, 2831, 0, 0, 0, 0, 1, 1),
		(drawing, 2830, 2830, 0, 0, 0, 0, 1, 1),
		(drawing, 2829, 2829, 0, 0, 0, 0, 1, 1),
		(drawing, 2828, 2828, 0, 0, 0, 0, 1, 1),
		(drawing, 2827, 2827, 0, 0, 0, 0, 1, 1),
		(drawing, 2826, 2826, 0, 0, 0, 0, 1, 1),
		(drawing, 2825, 2825, 0, 0, 0, 0, 1, 1),
		(drawing, 2824, 2824, 0, 0, 0, 0, 1, 1),
		(drawing, 2823, 2823, 0, 0, 0, 0, 1, 1),
		(drawing, 2822, 2822, 0, 0, 0, 0, 1, 1),
		(drawing, 2821, 2821, 0, 0, 0, 0, 1, 1),
		(drawing, 2820, 2820, 0, 0, 0, 0, 1, 1),
		(drawing, 2819, 2819, 0, 0, 0, 0, 1, 1),
		(drawing, 2818, 2818, 0, 0, 0, 0, 1, 1),
		(drawing, 2817, 2817, 0, 0, 0, 0, 1, 1),
		(drawing, 2816, 2816, 0, 0, 0, 0, 1, 1),
		(drawing, 2815, 2815, 0, 0, 0, 0, 1, 1),
		(drawing, 2814, 2814, 0, 0, 0, 0, 1, 1),
		(drawing, 2813, 2813, 0, 0, 0, 0, 1, 1),
		(drawing, 2812, 2812, 0, 0, 0, 0, 1, 1),
		(drawing, 2811, 2811, 0, 0, 0, 0, 1, 1),
		(drawing, 2810, 2810, 0, 0, 0, 0, 1, 1),
		(drawing, 2809, 2809, 0, 0, 0, 0, 1, 1),
		(drawing, 2808, 2808, 0, 0, 0, 0, 1, 1),
		(drawing, 2807, 2807, 0, 0, 0, 0, 1, 1),
		(drawing, 2806, 2806, 0, 0, 0, 0, 1, 1),
		(drawing, 2805, 2805, 0, 0, 0, 0, 1, 1),
		(drawing, 2804, 2804, 0, 0, 0, 0, 1, 1),
		(drawing, 2803, 2803, 0, 0, 0, 0, 1, 1),
		(drawing, 2802, 2802, 0, 0, 0, 0, 1, 1),
		(drawing, 2801, 2801, 0, 0, 0, 0, 1, 1),
		(drawing, 2800, 2800, 0, 0, 0, 0, 1, 1),
		(drawing, 2799, 2799, 0, 0, 0, 0, 1, 1),
		(drawing, 2798, 2798, 0, 0, 0, 0, 1, 1),
		(drawing, 2797, 2797, 0, 0, 0, 0, 1, 1),
		(drawing, 2796, 2796, 0, 0, 0, 0, 1, 1),
		(drawing, 2795, 2795, 0, 0, 0, 0, 1, 1),
		(drawing, 2794, 2794, 0, 0, 0, 0, 1, 1),
		(drawing, 2793, 2793, 0, 0, 0, 0, 1, 1),
		(drawing, 2792, 2792, 0, 0, 0, 0, 1, 1),
		(drawing, 2791, 2791, 0, 0, 0, 0, 1, 1),
		(drawing, 2790, 2790, 0, 0, 0, 0, 1, 1),
		(drawing, 2789, 2789, 0, 0, 0, 0, 1, 1),
		(drawing, 2788, 2788, 0, 0, 0, 0, 1, 1),
		(drawing, 2787, 2787, 0, 0, 0, 0, 1, 1),
		(drawing, 2786, 2786, 0, 0, 0, 0, 1, 1),
		(drawing, 2785, 2785, 0, 0, 0, 0, 1, 1),
		(drawing, 2784, 2784, 0, 0, 0, 0, 1, 1),
		(drawing, 2783, 2783, 0, 0, 0, 0, 1, 1),
		(drawing, 2782, 2782, 0, 0, 0, 0, 1, 1),
		(drawing, 2781, 2781, 0, 0, 0, 0, 1, 1),
		(drawing, 2780, 2780, 0, 0, 0, 0, 1, 1),
		(drawing, 2779, 2779, 0, 0, 0, 0, 1, 1),
		(drawing, 2778, 2778, 0, 0, 0, 0, 1, 1),
		(drawing, 2777, 2777, 0, 0, 0, 0, 1, 1),
		(drawing, 2776, 2776, 0, 0, 0, 0, 1, 1),
		(drawing, 2775, 2775, 0, 0, 0, 0, 1, 1),
		(drawing, 2774, 2774, 0, 0, 0, 0, 1, 1),
		(drawing, 2773, 2773, 0, 0, 0, 0, 1, 1),
		(drawing, 2772, 2772, 0, 0, 0, 0, 1, 1),
		(drawing, 2771, 2771, 0, 0, 0, 0, 1, 1),
		(drawing, 2770, 2770, 0, 0, 0, 0, 1, 1),
		(drawing, 2769, 2769, 0, 0, 0, 0, 1, 1),
		(drawing, 2768, 2768, 0, 0, 0, 0, 1, 1),
		(drawing, 2767, 2767, 0, 0, 0, 0, 1, 1),
		(drawing, 2766, 2766, 0, 0, 0, 0, 1, 1),
		(drawing, 2765, 2765, 0, 0, 0, 0, 1, 1),
		(drawing, 2764, 2764, 0, 0, 0, 0, 1, 1),
		(drawing, 2763, 2763, 0, 0, 0, 0, 1, 1),
		(drawing, 2762, 2762, 0, 0, 0, 0, 1, 1),
		(drawing, 2761, 2761, 0, 0, 0, 0, 1, 1),
		(drawing, 2760, 2760, 0, 0, 0, 0, 1, 1),
		(drawing, 2759, 2759, 0, 0, 0, 0, 1, 1),
		(drawing, 2758, 2758, 0, 0, 0, 0, 1, 1),
		(drawing, 2757, 2757, 0, 0, 0, 0, 1, 1),
		(drawing, 2756, 2756, 0, 0, 0, 0, 1, 1),
		(drawing, 2755, 2755, 0, 0, 0, 0, 1, 1),
		(drawing, 2754, 2754, 0, 0, 0, 0, 1, 1),
		(drawing, 2753, 2753, 0, 0, 0, 0, 1, 1),
		(drawing, 2752, 2752, 0, 0, 0, 0, 1, 1),
		(drawing, 2751, 2751, 0, 0, 0, 0, 1, 1),
		(drawing, 2750, 2750, 0, 0, 0, 0, 1, 1),
		(drawing, 2749, 2749, 0, 0, 0, 0, 1, 1),
		(drawing, 2748, 2748, 0, 0, 0, 0, 1, 1),
		(drawing, 2747, 2747, 0, 0, 0, 0, 1, 1),
		(drawing, 2746, 2746, 0, 0, 0, 0, 1, 1),
		(drawing, 2745, 2745, 0, 0, 0, 0, 1, 1),
		(drawing, 2744, 2744, 0, 0, 0, 0, 1, 1),
		(drawing, 2743, 2743, 0, 0, 0, 0, 1, 1),
		(drawing, 2742, 2742, 0, 0, 0, 0, 1, 1),
		(drawing, 2741, 2741, 0, 0, 0, 0, 1, 1),
		(drawing, 2740, 2740, 0, 0, 0, 0, 1, 1),
		(drawing, 2739, 2739, 0, 0, 0, 0, 1, 1),
		(drawing, 2738, 2738, 0, 0, 0, 0, 1, 1),
		(drawing, 2737, 2737, 0, 0, 0, 0, 1, 1),
		(drawing, 2736, 2736, 0, 0, 0, 0, 1, 1),
		(drawing, 2735, 2735, 0, 0, 0, 0, 1, 1),
		(drawing, 2734, 2734, 0, 0, 0, 0, 1, 1),
		(drawing, 2733, 2733, 0, 0, 0, 0, 1, 1),
		(drawing, 2732, 2732, 0, 0, 0, 0, 1, 1),
		(drawing, 2731, 2731, 0, 0, 0, 0, 1, 1),
		(drawing, 2730, 2730, 0, 0, 0, 0, 1, 1),
		(drawing, 2729, 2729, 0, 0, 0, 0, 1, 1),
		(drawing, 2728, 2728, 0, 0, 0, 0, 1, 1),
		(drawing, 2727, 2727, 0, 0, 0, 0, 1, 1),
		(drawing, 2726, 2726, 0, 0, 0, 0, 1, 1),
		(drawing, 2725, 2725, 0, 0, 0, 0, 1, 1),
		(drawing, 2724, 2724, 0, 0, 0, 0, 1, 1),
		(drawing, 2723, 2723, 0, 0, 0, 0, 1, 1),
		(drawing, 2722, 2722, 0, 0, 0, 0, 1, 1),
		(drawing, 2721, 2721, 0, 0, 0, 0, 1, 1),
		(drawing, 2720, 2720, 0, 0, 0, 0, 1, 1),
		(drawing, 2719, 2719, 0, 0, 0, 0, 1, 1),
		(drawing, 2718, 2718, 0, 0, 0, 0, 1, 1),
		(drawing, 2717, 2717, 0, 0, 0, 0, 1, 1),
		(drawing, 2716, 2716, 0, 0, 0, 0, 1, 1),
		(drawing, 2715, 2715, 0, 0, 0, 0, 1, 1),
		(drawing, 2714, 2714, 0, 0, 0, 0, 1, 1),
		(drawing, 2713, 2713, 0, 0, 0, 0, 1, 1),
		(drawing, 2712, 2712, 0, 0, 0, 0, 1, 1),
		(drawing, 2711, 2711, 0, 0, 0, 0, 1, 1),
		(drawing, 2710, 2710, 0, 0, 0, 0, 1, 1),
		(drawing, 2709, 2709, 0, 0, 0, 0, 1, 1),
		(drawing, 2708, 2708, 0, 0, 0, 0, 1, 1),
		(drawing, 2707, 2707, 0, 0, 0, 0, 1, 1),
		(drawing, 2706, 2706, 0, 0, 0, 0, 1, 1),
		(drawing, 2705, 2705, 0, 0, 0, 0, 1, 1),
		(drawing, 2704, 2704, 0, 0, 0, 0, 1, 1),
		(drawing, 2703, 2703, 0, 0, 0, 0, 1, 1),
		(drawing, 2702, 2702, 0, 0, 0, 0, 1, 1),
		(drawing, 2701, 2701, 0, 0, 0, 0, 1, 1),
		(drawing, 2700, 2700, 0, 0, 0, 0, 1, 1),
		(drawing, 2699, 2699, 0, 0, 0, 0, 1, 1),
		(drawing, 2698, 2698, 0, 0, 0, 0, 1, 1),
		(drawing, 2697, 2697, 0, 0, 0, 0, 1, 1),
		(drawing, 2696, 2696, 0, 0, 0, 0, 1, 1),
		(drawing, 2695, 2695, 0, 0, 0, 0, 1, 1),
		(drawing, 2694, 2694, 0, 0, 0, 0, 1, 1),
		(drawing, 2693, 2693, 0, 0, 0, 0, 1, 1),
		(drawing, 2692, 2692, 0, 0, 0, 0, 1, 1),
		(drawing, 2691, 2691, 0, 0, 0, 0, 1, 1),
		(drawing, 2690, 2690, 0, 0, 0, 0, 1, 1),
		(drawing, 2689, 2689, 0, 0, 0, 0, 1, 1),
		(drawing, 2688, 2688, 0, 0, 0, 0, 1, 1),
		(drawing, 2687, 2687, 0, 0, 0, 0, 1, 1),
		(drawing, 2686, 2686, 0, 0, 0, 0, 1, 1),
		(drawing, 2685, 2685, 0, 0, 0, 0, 1, 1),
		(drawing, 2684, 2684, 0, 0, 0, 0, 1, 1),
		(drawing, 2683, 2683, 0, 0, 0, 0, 1, 1),
		(drawing, 2682, 2682, 0, 0, 0, 0, 1, 1),
		(drawing, 2681, 2681, 0, 0, 0, 0, 1, 1),
		(drawing, 2680, 2680, 0, 0, 0, 0, 1, 1),
		(drawing, 2679, 2679, 0, 0, 0, 0, 1, 1),
		(drawing, 2678, 2678, 0, 0, 0, 0, 1, 1),
		(drawing, 2677, 2677, 0, 0, 0, 0, 1, 1),
		(drawing, 2676, 2676, 0, 0, 0, 0, 1, 1),
		(drawing, 2675, 2675, 0, 0, 0, 0, 1, 1),
		(drawing, 2674, 2674, 0, 0, 0, 0, 1, 1),
		(drawing, 2673, 2673, 0, 0, 0, 0, 1, 1),
		(drawing, 2672, 2672, 0, 0, 0, 0, 1, 1),
		(drawing, 2671, 2671, 0, 0, 0, 0, 1, 1),
		(drawing, 2670, 2670, 0, 0, 0, 0, 1, 1),
		(drawing, 2669, 2669, 0, 0, 0, 0, 1, 1),
		(drawing, 2668, 2668, 0, 0, 0, 0, 1, 1),
		(drawing, 2667, 2667, 0, 0, 0, 0, 1, 1),
		(drawing, 2666, 2666, 0, 0, 0, 0, 1, 1),
		(drawing, 2665, 2665, 0, 0, 0, 0, 1, 1),
		(drawing, 2664, 2664, 0, 0, 0, 0, 1, 1),
		(drawing, 2663, 2663, 0, 0, 0, 0, 1, 1),
		(drawing, 2662, 2662, 0, 0, 0, 0, 1, 1),
		(drawing, 2661, 2661, 0, 0, 0, 0, 1, 1),
		(drawing, 2660, 2660, 0, 0, 0, 0, 1, 1),
		(drawing, 2659, 2659, 0, 0, 0, 0, 1, 1),
		(drawing, 2658, 2658, 0, 0, 0, 0, 1, 1),
		(drawing, 2657, 2657, 0, 0, 0, 0, 1, 1),
		(drawing, 2656, 2656, 0, 0, 0, 0, 1, 1),
		(drawing, 2655, 2655, 0, 0, 0, 0, 1, 1),
		(drawing, 2654, 2654, 0, 0, 0, 0, 1, 1),
		(drawing, 2653, 2653, 0, 0, 0, 0, 1, 1),
		(drawing, 2652, 2652, 0, 0, 0, 0, 1, 1),
		(drawing, 2651, 2651, 0, 0, 0, 0, 1, 1),
		(drawing, 2650, 2650, 0, 0, 0, 0, 1, 1),
		(drawing, 2649, 2649, 0, 0, 0, 0, 1, 1),
		(drawing, 2648, 2648, 0, 0, 0, 0, 1, 1),
		(drawing, 2647, 2647, 0, 0, 0, 0, 1, 1),
		(drawing, 2646, 2646, 0, 0, 0, 0, 1, 1),
		(drawing, 2645, 2645, 0, 0, 0, 0, 1, 1),
		(drawing, 2644, 2644, 0, 0, 0, 0, 1, 1),
		(drawing, 2643, 2643, 0, 0, 0, 0, 1, 1),
		(drawing, 2642, 2642, 0, 0, 0, 0, 1, 1),
		(drawing, 2641, 2641, 0, 0, 0, 0, 1, 1),
		(drawing, 2640, 2640, 0, 0, 0, 0, 1, 1),
		(drawing, 2639, 2639, 0, 0, 0, 0, 1, 1),
		(drawing, 2638, 2638, 0, 0, 0, 0, 1, 1),
		(drawing, 2637, 2637, 0, 0, 0, 0, 1, 1),
		(drawing, 2636, 2636, 0, 0, 0, 0, 1, 1),
		(drawing, 2635, 2635, 0, 0, 0, 0, 1, 1),
		(drawing, 2634, 2634, 0, 0, 0, 0, 1, 1),
		(drawing, 2633, 2633, 0, 0, 0, 0, 1, 1),
		(drawing, 2632, 2632, 0, 0, 0, 0, 1, 1),
		(drawing, 2631, 2631, 0, 0, 0, 0, 1, 1),
		(drawing, 2630, 2630, 0, 0, 0, 0, 1, 1),
		(drawing, 2629, 2629, 0, 0, 0, 0, 1, 1),
		(drawing, 2628, 2628, 0, 0, 0, 0, 1, 1),
		(drawing, 2627, 2627, 0, 0, 0, 0, 1, 1),
		(drawing, 2626, 2626, 0, 0, 0, 0, 1, 1),
		(drawing, 2625, 2625, 0, 0, 0, 0, 1, 1),
		(drawing, 2624, 2624, 0, 0, 0, 0, 1, 1),
		(drawing, 2623, 2623, 0, 0, 0, 0, 1, 1),
		(drawing, 2622, 2622, 0, 0, 0, 0, 1, 1),
		(drawing, 2621, 2621, 0, 0, 0, 0, 1, 1),
		(drawing, 2620, 2620, 0, 0, 0, 0, 1, 1),
		(drawing, 2619, 2619, 0, 0, 0, 0, 1, 1),
		(drawing, 2618, 2618, 0, 0, 0, 0, 1, 1),
		(drawing, 2617, 2617, 0, 0, 0, 0, 1, 1),
		(drawing, 2616, 2616, 0, 0, 0, 0, 1, 1),
		(drawing, 2615, 2615, 0, 0, 0, 0, 1, 1),
		(drawing, 2614, 2614, 0, 0, 0, 0, 1, 1),
		(drawing, 2613, 2613, 0, 0, 0, 0, 1, 1),
		(drawing, 2612, 2612, 0, 0, 0, 0, 1, 1),
		(drawing, 2611, 2611, 0, 0, 0, 0, 1, 1),
		(drawing, 2610, 2610, 0, 0, 0, 0, 1, 1),
		(drawing, 2609, 2609, 0, 0, 0, 0, 1, 1),
		(drawing, 2608, 2608, 0, 0, 0, 0, 1, 1),
		(drawing, 2607, 2607, 0, 0, 0, 0, 1, 1),
		(drawing, 2606, 2606, 0, 0, 0, 0, 1, 1),
		(drawing, 2605, 2605, 0, 0, 0, 0, 1, 1),
		(drawing, 2604, 2604, 0, 0, 0, 0, 1, 1),
		(drawing, 2603, 2603, 0, 0, 0, 0, 1, 1),
		(drawing, 2602, 2602, 0, 0, 0, 0, 1, 1),
		(drawing, 2601, 2601, 0, 0, 0, 0, 1, 1),
		(drawing, 2600, 2600, 0, 0, 0, 0, 1, 1),
		(drawing, 2599, 2599, 0, 0, 0, 0, 1, 1),
		(drawing, 2598, 2598, 0, 0, 0, 0, 1, 1),
		(drawing, 2597, 2597, 0, 0, 0, 0, 1, 1),
		(drawing, 2596, 2596, 0, 0, 0, 0, 1, 1),
		(drawing, 2595, 2595, 0, 0, 0, 0, 1, 1),
		(drawing, 2594, 2594, 0, 0, 0, 0, 1, 1),
		(drawing, 2593, 2593, 0, 0, 0, 0, 1, 1),
		(drawing, 2592, 2592, 0, 0, 0, 0, 1, 1),
		(drawing, 2591, 2591, 0, 0, 0, 0, 1, 1),
		(drawing, 2590, 2590, 0, 0, 0, 0, 1, 1),
		(drawing, 2589, 2589, 0, 0, 0, 0, 1, 1),
		(drawing, 2588, 2588, 0, 0, 0, 0, 1, 1),
		(drawing, 2587, 2587, 0, 0, 0, 0, 1, 1),
		(drawing, 2586, 2586, 0, 0, 0, 0, 1, 1),
		(drawing, 2585, 2585, 0, 0, 0, 0, 1, 1),
		(drawing, 2584, 2584, 0, 0, 0, 0, 1, 1),
		(drawing, 2583, 2583, 0, 0, 0, 0, 1, 1),
		(drawing, 2582, 2582, 0, 0, 0, 0, 1, 1),
		(drawing, 2581, 2581, 0, 0, 0, 0, 1, 1),
		(drawing, 2580, 2580, 0, 0, 0, 0, 1, 1),
		(drawing, 2579, 2579, 0, 0, 0, 0, 1, 1),
		(drawing, 2578, 2578, 0, 0, 0, 0, 1, 1),
		(drawing, 2577, 2577, 0, 0, 0, 0, 1, 1),
		(drawing, 2576, 2576, 0, 0, 0, 0, 1, 1),
		(drawing, 2575, 2575, 0, 0, 0, 0, 1, 1),
		(drawing, 2574, 2574, 0, 0, 0, 0, 1, 1),
		(drawing, 2573, 2573, 0, 0, 0, 0, 1, 1),
		(drawing, 2572, 2572, 0, 0, 0, 0, 1, 1),
		(drawing, 2571, 2571, 0, 0, 0, 0, 1, 1),
		(drawing, 2570, 2570, 0, 0, 0, 0, 1, 1),
		(drawing, 2569, 2569, 0, 0, 0, 0, 1, 1),
		(drawing, 2568, 2568, 0, 0, 0, 0, 1, 1),
		(drawing, 2567, 2567, 0, 0, 0, 0, 1, 1),
		(drawing, 2566, 2566, 0, 0, 0, 0, 1, 1),
		(drawing, 2565, 2565, 0, 0, 0, 0, 1, 1),
		(drawing, 2564, 2564, 0, 0, 0, 0, 1, 1),
		(drawing, 2563, 2563, 0, 0, 0, 0, 1, 1),
		(drawing, 2562, 2562, 0, 0, 0, 0, 1, 1),
		(drawing, 2561, 2561, 0, 0, 0, 0, 1, 1),
		(drawing, 2560, 2560, 0, 0, 0, 0, 1, 1),
		(drawing, 2559, 2559, 0, 0, 0, 0, 1, 1),
		(drawing, 2558, 2558, 0, 0, 0, 0, 1, 1),
		(drawing, 2557, 2557, 0, 0, 0, 0, 1, 1),
		(drawing, 2556, 2556, 0, 0, 0, 0, 1, 1),
		(drawing, 2555, 2555, 0, 0, 0, 0, 1, 1),
		(drawing, 2554, 2554, 0, 0, 0, 0, 1, 1),
		(drawing, 2553, 2553, 0, 0, 0, 0, 1, 1),
		(drawing, 2552, 2552, 0, 0, 0, 0, 1, 1),
		(drawing, 2551, 2551, 0, 0, 0, 0, 1, 1),
		(drawing, 2550, 2550, 0, 0, 0, 0, 1, 1),
		(drawing, 2549, 2549, 0, 0, 0, 0, 1, 1),
		(drawing, 2548, 2548, 0, 0, 0, 0, 1, 1),
		(drawing, 2547, 2547, 0, 0, 0, 0, 1, 1),
		(drawing, 2546, 2546, 0, 0, 0, 0, 1, 1),
		(drawing, 2545, 2545, 0, 0, 0, 0, 1, 1),
		(drawing, 2544, 2544, 0, 0, 0, 0, 1, 1),
		(drawing, 2543, 2543, 0, 0, 0, 0, 1, 1),
		(drawing, 2542, 2542, 0, 0, 0, 0, 1, 1),
		(drawing, 2541, 2541, 0, 0, 0, 0, 1, 1),
		(drawing, 2540, 2540, 0, 0, 0, 0, 1, 1),
		(drawing, 2539, 2539, 0, 0, 0, 0, 1, 1),
		(drawing, 2538, 2538, 0, 0, 0, 0, 1, 1),
		(drawing, 2537, 2537, 0, 0, 0, 0, 1, 1),
		(drawing, 2536, 2536, 0, 0, 0, 0, 1, 1),
		(drawing, 2535, 2535, 0, 0, 0, 0, 1, 1),
		(drawing, 2534, 2534, 0, 0, 0, 0, 1, 1),
		(drawing, 2533, 2533, 0, 0, 0, 0, 1, 1),
		(drawing, 2532, 2532, 0, 0, 0, 0, 1, 1),
		(drawing, 2531, 2531, 0, 0, 0, 0, 1, 1),
		(drawing, 2530, 2530, 0, 0, 0, 0, 1, 1),
		(drawing, 2529, 2529, 0, 0, 0, 0, 1, 1),
		(drawing, 2528, 2528, 0, 0, 0, 0, 1, 1),
		(drawing, 2527, 2527, 0, 0, 0, 0, 1, 1),
		(drawing, 2526, 2526, 0, 0, 0, 0, 1, 1),
		(drawing, 2525, 2525, 0, 0, 0, 0, 1, 1),
		(drawing, 2524, 2524, 0, 0, 0, 0, 1, 1),
		(drawing, 2523, 2523, 0, 0, 0, 0, 1, 1),
		(drawing, 2522, 2522, 0, 0, 0, 0, 1, 1),
		(drawing, 2521, 2521, 0, 0, 0, 0, 1, 1),
		(drawing, 2520, 2520, 0, 0, 0, 0, 1, 1),
		(drawing, 2519, 2519, 0, 0, 0, 0, 1, 1),
		(drawing, 2518, 2518, 0, 0, 0, 0, 1, 1),
		(drawing, 2517, 2517, 0, 0, 0, 0, 1, 1),
		(drawing, 2516, 2516, 0, 0, 0, 0, 1, 1),
		(drawing, 2515, 2515, 0, 0, 0, 0, 1, 1),
		(drawing, 2514, 2514, 0, 0, 0, 0, 1, 1),
		(drawing, 2513, 2513, 0, 0, 0, 0, 1, 1),
		(drawing, 2512, 2512, 0, 0, 0, 0, 1, 1),
		(drawing, 2511, 2511, 0, 0, 0, 0, 1, 1),
		(drawing, 2510, 2510, 0, 0, 0, 0, 1, 1),
		(drawing, 2509, 2509, 0, 0, 0, 0, 1, 1),
		(drawing, 2508, 2508, 0, 0, 0, 0, 1, 1),
		(drawing, 2507, 2507, 0, 0, 0, 0, 1, 1),
		(drawing, 2506, 2506, 0, 0, 0, 0, 1, 1),
		(drawing, 2505, 2505, 0, 0, 0, 0, 1, 1),
		(drawing, 2504, 2504, 0, 0, 0, 0, 1, 1),
		(drawing, 2503, 2503, 0, 0, 0, 0, 1, 1),
		(drawing, 2502, 2502, 0, 0, 0, 0, 1, 1),
		(drawing, 2501, 2501, 0, 0, 0, 0, 1, 1),
		(drawing, 2500, 2500, 0, 0, 0, 0, 1, 1),
		(drawing, 2499, 2499, 0, 0, 0, 0, 1, 1),
		(drawing, 2498, 2498, 0, 0, 0, 0, 1, 1),
		(drawing, 2497, 2497, 0, 0, 0, 0, 1, 1),
		(drawing, 2496, 2496, 0, 0, 0, 0, 1, 1),
		(drawing, 2495, 2495, 0, 0, 0, 0, 1, 1),
		(drawing, 2494, 2494, 0, 0, 0, 0, 1, 1),
		(drawing, 2493, 2493, 0, 0, 0, 0, 1, 1),
		(drawing, 2492, 2492, 0, 0, 0, 0, 1, 1),
		(drawing, 2491, 2491, 0, 0, 0, 0, 1, 1),
		(drawing, 2490, 2490, 0, 0, 0, 0, 1, 1),
		(drawing, 2489, 2489, 0, 0, 0, 0, 1, 1),
		(drawing, 2488, 2488, 0, 0, 0, 0, 1, 1),
		(drawing, 2487, 2487, 0, 0, 0, 0, 1, 1),
		(drawing, 2486, 2486, 0, 0, 0, 0, 1, 1),
		(drawing, 2485, 2485, 0, 0, 0, 0, 1, 1),
		(drawing, 2484, 2484, 0, 0, 0, 0, 1, 1),
		(drawing, 2483, 2483, 0, 0, 0, 0, 1, 1),
		(drawing, 2482, 2482, 0, 0, 0, 0, 1, 1),
		(drawing, 2481, 2481, 0, 0, 0, 0, 1, 1),
		(drawing, 2480, 2480, 0, 0, 0, 0, 1, 1),
		(drawing, 2479, 2479, 0, 0, 0, 0, 1, 1),
		(drawing, 2478, 2478, 0, 0, 0, 0, 1, 1),
		(drawing, 2477, 2477, 0, 0, 0, 0, 1, 1),
		(drawing, 2476, 2476, 0, 0, 0, 0, 1, 1),
		(drawing, 2475, 2475, 0, 0, 0, 0, 1, 1),
		(drawing, 2474, 2474, 0, 0, 0, 0, 1, 1),
		(drawing, 2473, 2473, 0, 0, 0, 0, 1, 1),
		(drawing, 2472, 2472, 0, 0, 0, 0, 1, 1),
		(drawing, 2471, 2471, 0, 0, 0, 0, 1, 1),
		(drawing, 2470, 2470, 0, 0, 0, 0, 1, 1),
		(drawing, 2469, 2469, 0, 0, 0, 0, 1, 1),
		(drawing, 2468, 2468, 0, 0, 0, 0, 1, 1),
		(drawing, 2467, 2467, 0, 0, 0, 0, 1, 1),
		(drawing, 2466, 2466, 0, 0, 0, 0, 1, 1),
		(drawing, 2465, 2465, 0, 0, 0, 0, 1, 1),
		(drawing, 2464, 2464, 0, 0, 0, 0, 1, 1),
		(drawing, 2463, 2463, 0, 0, 0, 0, 1, 1),
		(drawing, 2462, 2462, 0, 0, 0, 0, 1, 1),
		(drawing, 2461, 2461, 0, 0, 0, 0, 1, 1),
		(drawing, 2460, 2460, 0, 0, 0, 0, 1, 1),
		(drawing, 2459, 2459, 0, 0, 0, 0, 1, 1),
		(drawing, 2458, 2458, 0, 0, 0, 0, 1, 1),
		(drawing, 2457, 2457, 0, 0, 0, 0, 1, 1),
		(drawing, 2456, 2456, 0, 0, 0, 0, 1, 1),
		(drawing, 2455, 2455, 0, 0, 0, 0, 1, 1),
		(drawing, 2454, 2454, 0, 0, 0, 0, 1, 1),
		(drawing, 2453, 2453, 0, 0, 0, 0, 1, 1),
		(drawing, 2452, 2452, 0, 0, 0, 0, 1, 1),
		(drawing, 2451, 2451, 0, 0, 0, 0, 1, 1),
		(drawing, 2450, 2450, 0, 0, 0, 0, 1, 1),
		(drawing, 2449, 2449, 0, 0, 0, 0, 1, 1),
		(drawing, 2448, 2448, 0, 0, 0, 0, 1, 1),
		(drawing, 2447, 2447, 0, 0, 0, 0, 1, 1),
		(drawing, 2446, 2446, 0, 0, 0, 0, 1, 1),
		(drawing, 2445, 2445, 0, 0, 0, 0, 1, 1),
		(drawing, 2444, 2444, 0, 0, 0, 0, 1, 1),
		(drawing, 2443, 2443, 0, 0, 0, 0, 1, 1),
		(drawing, 2442, 2442, 0, 0, 0, 0, 1, 1),
		(drawing, 2441, 2441, 0, 0, 0, 0, 1, 1),
		(drawing, 2440, 2440, 0, 0, 0, 0, 1, 1),
		(drawing, 2439, 2439, 0, 0, 0, 0, 1, 1),
		(drawing, 2438, 2438, 0, 0, 0, 0, 1, 1),
		(drawing, 2437, 2437, 0, 0, 0, 0, 1, 1),
		(drawing, 2436, 2436, 0, 0, 0, 0, 1, 1),
		(drawing, 2435, 2435, 0, 0, 0, 0, 1, 1),
		(drawing, 2434, 2434, 0, 0, 0, 0, 1, 1),
		(drawing, 2433, 2433, 0, 0, 0, 0, 1, 1),
		(drawing, 2432, 2432, 0, 0, 0, 0, 1, 1),
		(drawing, 2431, 2431, 0, 0, 0, 0, 1, 1),
		(drawing, 2430, 2430, 0, 0, 0, 0, 1, 1),
		(drawing, 2429, 2429, 0, 0, 0, 0, 1, 1),
		(drawing, 2428, 2428, 0, 0, 0, 0, 1, 1),
		(drawing, 2427, 2427, 0, 0, 0, 0, 1, 1),
		(drawing, 2426, 2426, 0, 0, 0, 0, 1, 1),
		(drawing, 2425, 2425, 0, 0, 0, 0, 1, 1),
		(drawing, 2424, 2424, 0, 0, 0, 0, 1, 1),
		(drawing, 2423, 2423, 0, 0, 0, 0, 1, 1),
		(drawing, 2422, 2422, 0, 0, 0, 0, 1, 1),
		(drawing, 2421, 2421, 0, 0, 0, 0, 1, 1),
		(drawing, 2420, 2420, 0, 0, 0, 0, 1, 1),
		(drawing, 2419, 2419, 0, 0, 0, 0, 1, 1),
		(drawing, 2418, 2418, 0, 0, 0, 0, 1, 1),
		(drawing, 2417, 2417, 0, 0, 0, 0, 1, 1),
		(drawing, 2416, 2416, 0, 0, 0, 0, 1, 1),
		(drawing, 2415, 2415, 0, 0, 0, 0, 1, 1),
		(drawing, 2414, 2414, 0, 0, 0, 0, 1, 1),
		(drawing, 2413, 2413, 0, 0, 0, 0, 1, 1),
		(drawing, 2412, 2412, 0, 0, 0, 0, 1, 1),
		(drawing, 2411, 2411, 0, 0, 0, 0, 1, 1),
		(drawing, 2410, 2410, 0, 0, 0, 0, 1, 1),
		(drawing, 2409, 2409, 0, 0, 0, 0, 1, 1),
		(drawing, 2408, 2408, 0, 0, 0, 0, 1, 1),
		(drawing, 2407, 2407, 0, 0, 0, 0, 1, 1),
		(drawing, 2406, 2406, 0, 0, 0, 0, 1, 1),
		(drawing, 2405, 2405, 0, 0, 0, 0, 1, 1),
		(drawing, 2404, 2404, 0, 0, 0, 0, 1, 1),
		(drawing, 2403, 2403, 0, 0, 0, 0, 1, 1),
		(drawing, 2402, 2402, 0, 0, 0, 0, 1, 1),
		(drawing, 2401, 2401, 0, 0, 0, 0, 1, 1),
		(drawing, 2400, 2400, 0, 0, 0, 0, 1, 1),
		(drawing, 2399, 2399, 0, 0, 0, 0, 1, 1),
		(drawing, 2398, 2398, 0, 0, 0, 0, 1, 1),
		(drawing, 2397, 2397, 0, 0, 0, 0, 1, 1),
		(drawing, 2396, 2396, 0, 0, 0, 0, 1, 1),
		(drawing, 2395, 2395, 0, 0, 0, 0, 1, 1),
		(drawing, 2394, 2394, 0, 0, 0, 0, 1, 1),
		(drawing, 2393, 2393, 0, 0, 0, 0, 1, 1),
		(drawing, 2392, 2392, 0, 0, 0, 0, 1, 1),
		(drawing, 2391, 2391, 0, 0, 0, 0, 1, 1),
		(drawing, 2390, 2390, 0, 0, 0, 0, 1, 1),
		(drawing, 2389, 2389, 0, 0, 0, 0, 1, 1),
		(drawing, 2388, 2388, 0, 0, 0, 0, 1, 1),
		(drawing, 2387, 2387, 0, 0, 0, 0, 1, 1),
		(drawing, 2386, 2386, 0, 0, 0, 0, 1, 1),
		(drawing, 2385, 2385, 0, 0, 0, 0, 1, 1),
		(drawing, 2384, 2384, 0, 0, 0, 0, 1, 1),
		(drawing, 2383, 2383, 0, 0, 0, 0, 1, 1),
		(drawing, 2382, 2382, 0, 0, 0, 0, 1, 1),
		(drawing, 2381, 2381, 0, 0, 0, 0, 1, 1),
		(drawing, 2380, 2380, 0, 0, 0, 0, 1, 1),
		(drawing, 2379, 2379, 0, 0, 0, 0, 1, 1),
		(drawing, 2378, 2378, 0, 0, 0, 0, 1, 1),
		(drawing, 2377, 2377, 0, 0, 0, 0, 1, 1),
		(drawing, 2376, 2376, 0, 0, 0, 0, 1, 1),
		(drawing, 2375, 2375, 0, 0, 0, 0, 1, 1),
		(drawing, 2374, 2374, 0, 0, 0, 0, 1, 1),
		(drawing, 2373, 2373, 0, 0, 0, 0, 1, 1),
		(drawing, 2372, 2372, 0, 0, 0, 0, 1, 1),
		(drawing, 2371, 2371, 0, 0, 0, 0, 1, 1),
		(drawing, 2370, 2370, 0, 0, 0, 0, 1, 1),
		(drawing, 2369, 2369, 0, 0, 0, 0, 1, 1),
		(drawing, 2368, 2368, 0, 0, 0, 0, 1, 1),
		(drawing, 2367, 2367, 0, 0, 0, 0, 1, 1),
		(drawing, 2366, 2366, 0, 0, 0, 0, 1, 1),
		(drawing, 2365, 2365, 0, 0, 0, 0, 1, 1),
		(drawing, 2364, 2364, 0, 0, 0, 0, 1, 1),
		(drawing, 2363, 2363, 0, 0, 0, 0, 1, 1),
		(drawing, 2362, 2362, 0, 0, 0, 0, 1, 1),
		(drawing, 2361, 2361, 0, 0, 0, 0, 1, 1),
		(drawing, 2360, 2360, 0, 0, 0, 0, 1, 1),
		(drawing, 2359, 2359, 0, 0, 0, 0, 1, 1),
		(drawing, 2358, 2358, 0, 0, 0, 0, 1, 1),
		(drawing, 2357, 2357, 0, 0, 0, 0, 1, 1),
		(drawing, 2356, 2356, 0, 0, 0, 0, 1, 1),
		(drawing, 2355, 2355, 0, 0, 0, 0, 1, 1),
		(drawing, 2354, 2354, 0, 0, 0, 0, 1, 1),
		(drawing, 2353, 2353, 0, 0, 0, 0, 1, 1),
		(drawing, 2352, 2352, 0, 0, 0, 0, 1, 1),
		(drawing, 2351, 2351, 0, 0, 0, 0, 1, 1),
		(drawing, 2350, 2350, 0, 0, 0, 0, 1, 1),
		(drawing, 2349, 2349, 0, 0, 0, 0, 1, 1),
		(drawing, 2348, 2348, 0, 0, 0, 0, 1, 1),
		(drawing, 2347, 2347, 0, 0, 0, 0, 1, 1),
		(drawing, 2346, 2346, 0, 0, 0, 0, 1, 1),
		(drawing, 2345, 2345, 0, 0, 0, 0, 1, 1),
		(drawing, 2344, 2344, 0, 0, 0, 0, 1, 1),
		(drawing, 2343, 2343, 0, 0, 0, 0, 1, 1),
		(drawing, 2342, 2342, 0, 0, 0, 0, 1, 1),
		(drawing, 2341, 2341, 0, 0, 0, 0, 1, 1),
		(drawing, 2340, 2340, 0, 0, 0, 0, 1, 1),
		(drawing, 2339, 2339, 0, 0, 0, 0, 1, 1),
		(drawing, 2338, 2338, 0, 0, 0, 0, 1, 1),
		(drawing, 2337, 2337, 0, 0, 0, 0, 1, 1),
		(drawing, 2336, 2336, 0, 0, 0, 0, 1, 1),
		(drawing, 2335, 2335, 0, 0, 0, 0, 1, 1),
		(drawing, 2334, 2334, 0, 0, 0, 0, 1, 1),
		(drawing, 2333, 2333, 0, 0, 0, 0, 1, 1),
		(drawing, 2332, 2332, 0, 0, 0, 0, 1, 1),
		(drawing, 2331, 2331, 0, 0, 0, 0, 1, 1),
		(drawing, 2330, 2330, 0, 0, 0, 0, 1, 1),
		(drawing, 2329, 2329, 0, 0, 0, 0, 1, 1),
		(drawing, 2328, 2328, 0, 0, 0, 0, 1, 1),
		(drawing, 2327, 2327, 0, 0, 0, 0, 1, 1),
		(drawing, 2326, 2326, 0, 0, 0, 0, 1, 1),
		(drawing, 2325, 2325, 0, 0, 0, 0, 1, 1),
		(drawing, 2324, 2324, 0, 0, 0, 0, 1, 1),
		(drawing, 2323, 2323, 0, 0, 0, 0, 1, 1),
		(drawing, 2322, 2322, 0, 0, 0, 0, 1, 1),
		(drawing, 2321, 2321, 0, 0, 0, 0, 1, 1),
		(drawing, 2320, 2320, 0, 0, 0, 0, 1, 1),
		(drawing, 2319, 2319, 0, 0, 0, 0, 1, 1),
		(drawing, 2318, 2318, 0, 0, 0, 0, 1, 1),
		(drawing, 2317, 2317, 0, 0, 0, 0, 1, 1),
		(drawing, 2316, 2316, 0, 0, 0, 0, 1, 1),
		(drawing, 2315, 2315, 0, 0, 0, 0, 1, 1),
		(drawing, 2314, 2314, 0, 0, 0, 0, 1, 1),
		(drawing, 2313, 2313, 0, 0, 0, 0, 1, 1),
		(drawing, 2312, 2312, 0, 0, 0, 0, 1, 1),
		(drawing, 2311, 2311, 0, 0, 0, 0, 1, 1),
		(drawing, 2310, 2310, 0, 0, 0, 0, 1, 1),
		(drawing, 2309, 2309, 0, 0, 0, 0, 1, 1),
		(drawing, 2308, 2308, 0, 0, 0, 0, 1, 1),
		(drawing, 2307, 2307, 0, 0, 0, 0, 1, 1),
		(drawing, 2306, 2306, 0, 0, 0, 0, 1, 1),
		(drawing, 2305, 2305, 0, 0, 0, 0, 1, 1),
		(drawing, 2304, 2304, 0, 0, 0, 0, 1, 1),
		(drawing, 2303, 2303, 0, 0, 0, 0, 1, 1),
		(drawing, 2302, 2302, 0, 0, 0, 0, 1, 1),
		(drawing, 2301, 2301, 0, 0, 0, 0, 1, 1),
		(drawing, 2300, 2300, 0, 0, 0, 0, 1, 1),
		(drawing, 2299, 2299, 0, 0, 0, 0, 1, 1),
		(drawing, 2298, 2298, 0, 0, 0, 0, 1, 1),
		(drawing, 2297, 2297, 0, 0, 0, 0, 1, 1),
		(drawing, 2296, 2296, 0, 0, 0, 0, 1, 1),
		(drawing, 2295, 2295, 0, 0, 0, 0, 1, 1),
		(drawing, 2294, 2294, 0, 0, 0, 0, 1, 1),
		(drawing, 2293, 2293, 0, 0, 0, 0, 1, 1),
		(drawing, 2292, 2292, 0, 0, 0, 0, 1, 1),
		(drawing, 2291, 2291, 0, 0, 0, 0, 1, 1),
		(drawing, 2290, 2290, 0, 0, 0, 0, 1, 1),
		(drawing, 2289, 2289, 0, 0, 0, 0, 1, 1),
		(drawing, 2288, 2288, 0, 0, 0, 0, 1, 1),
		(drawing, 2287, 2287, 0, 0, 0, 0, 1, 1),
		(drawing, 2286, 2286, 0, 0, 0, 0, 1, 1),
		(drawing, 2285, 2285, 0, 0, 0, 0, 1, 1),
		(drawing, 2284, 2284, 0, 0, 0, 0, 1, 1),
		(drawing, 2283, 2283, 0, 0, 0, 0, 1, 1),
		(drawing, 2282, 2282, 0, 0, 0, 0, 1, 1),
		(drawing, 2281, 2281, 0, 0, 0, 0, 1, 1),
		(drawing, 2280, 2280, 0, 0, 0, 0, 1, 1),
		(drawing, 2279, 2279, 0, 0, 0, 0, 1, 1),
		(drawing, 2278, 2278, 0, 0, 0, 0, 1, 1),
		(drawing, 2277, 2277, 0, 0, 0, 0, 1, 1),
		(drawing, 2276, 2276, 0, 0, 0, 0, 1, 1),
		(drawing, 2275, 2275, 0, 0, 0, 0, 1, 1),
		(drawing, 2274, 2274, 0, 0, 0, 0, 1, 1),
		(drawing, 2273, 2273, 0, 0, 0, 0, 1, 1),
		(drawing, 2272, 2272, 0, 0, 0, 0, 1, 1),
		(drawing, 2271, 2271, 0, 0, 0, 0, 1, 1),
		(drawing, 2270, 2270, 0, 0, 0, 0, 1, 1),
		(drawing, 2269, 2269, 0, 0, 0, 0, 1, 1),
		(drawing, 2268, 2268, 0, 0, 0, 0, 1, 1),
		(drawing, 2267, 2267, 0, 0, 0, 0, 1, 1),
		(drawing, 2266, 2266, 0, 0, 0, 0, 1, 1),
		(drawing, 2265, 2265, 0, 0, 0, 0, 1, 1),
		(drawing, 2264, 2264, 0, 0, 0, 0, 1, 1),
		(drawing, 2263, 2263, 0, 0, 0, 0, 1, 1),
		(drawing, 2262, 2262, 0, 0, 0, 0, 1, 1),
		(drawing, 2261, 2261, 0, 0, 0, 0, 1, 1),
		(drawing, 2260, 2260, 0, 0, 0, 0, 1, 1),
		(drawing, 2259, 2259, 0, 0, 0, 0, 1, 1),
		(drawing, 2258, 2258, 0, 0, 0, 0, 1, 1),
		(drawing, 2257, 2257, 0, 0, 0, 0, 1, 1),
		(drawing, 2256, 2256, 0, 0, 0, 0, 1, 1),
		(drawing, 2255, 2255, 0, 0, 0, 0, 1, 1),
		(drawing, 2254, 2254, 0, 0, 0, 0, 1, 1),
		(drawing, 2253, 2253, 0, 0, 0, 0, 1, 1),
		(drawing, 2252, 2252, 0, 0, 0, 0, 1, 1),
		(drawing, 2251, 2251, 0, 0, 0, 0, 1, 1),
		(drawing, 2250, 2250, 0, 0, 0, 0, 1, 1),
		(drawing, 2249, 2249, 0, 0, 0, 0, 1, 1),
		(drawing, 2248, 2248, 0, 0, 0, 0, 1, 1),
		(drawing, 2247, 2247, 0, 0, 0, 0, 1, 1),
		(drawing, 2246, 2246, 0, 0, 0, 0, 1, 1),
		(drawing, 2245, 2245, 0, 0, 0, 0, 1, 1),
		(drawing, 2244, 2244, 0, 0, 0, 0, 1, 1),
		(drawing, 2243, 2243, 0, 0, 0, 0, 1, 1),
		(drawing, 2242, 2242, 0, 0, 0, 0, 1, 1),
		(drawing, 2241, 2241, 0, 0, 0, 0, 1, 1),
		(drawing, 2240, 2240, 0, 0, 0, 0, 1, 1),
		(drawing, 2239, 2239, 0, 0, 0, 0, 1, 1),
		(drawing, 2238, 2238, 0, 0, 0, 0, 1, 1),
		(drawing, 2237, 2237, 0, 0, 0, 0, 1, 1),
		(drawing, 2236, 2236, 0, 0, 0, 0, 1, 1),
		(drawing, 2235, 2235, 0, 0, 0, 0, 1, 1),
		(drawing, 2234, 2234, 0, 0, 0, 0, 1, 1),
		(drawing, 2233, 2233, 0, 0, 0, 0, 1, 1),
		(drawing, 2232, 2232, 0, 0, 0, 0, 1, 1),
		(drawing, 2231, 2231, 0, 0, 0, 0, 1, 1),
		(drawing, 2230, 2230, 0, 0, 0, 0, 1, 1),
		(drawing, 2229, 2229, 0, 0, 0, 0, 1, 1),
		(drawing, 2228, 2228, 0, 0, 0, 0, 1, 1),
		(drawing, 2227, 2227, 0, 0, 0, 0, 1, 1),
		(drawing, 2226, 2226, 0, 0, 0, 0, 1, 1),
		(drawing, 2225, 2225, 0, 0, 0, 0, 1, 1),
		(drawing, 2224, 2224, 0, 0, 0, 0, 1, 1),
		(drawing, 2223, 2223, 0, 0, 0, 0, 1, 1),
		(drawing, 2222, 2222, 0, 0, 0, 0, 1, 1),
		(drawing, 2221, 2221, 0, 0, 0, 0, 1, 1),
		(drawing, 2220, 2220, 0, 0, 0, 0, 1, 1),
		(drawing, 2219, 2219, 0, 0, 0, 0, 1, 1),
		(drawing, 2218, 2218, 0, 0, 0, 0, 1, 1),
		(drawing, 2217, 2217, 0, 0, 0, 0, 1, 1),
		(drawing, 2216, 2216, 0, 0, 0, 0, 1, 1),
		(drawing, 2215, 2215, 0, 0, 0, 0, 1, 1),
		(drawing, 2214, 2214, 0, 0, 0, 0, 1, 1),
		(drawing, 2213, 2213, 0, 0, 0, 0, 1, 1),
		(drawing, 2212, 2212, 0, 0, 0, 0, 1, 1),
		(drawing, 2211, 2211, 0, 0, 0, 0, 1, 1),
		(drawing, 2210, 2210, 0, 0, 0, 0, 1, 1),
		(drawing, 2209, 2209, 0, 0, 0, 0, 1, 1),
		(drawing, 2208, 2208, 0, 0, 0, 0, 1, 1),
		(drawing, 2207, 2207, 0, 0, 0, 0, 1, 1),
		(drawing, 2206, 2206, 0, 0, 0, 0, 1, 1),
		(drawing, 2205, 2205, 0, 0, 0, 0, 1, 1),
		(drawing, 2204, 2204, 0, 0, 0, 0, 1, 1),
		(drawing, 2203, 2203, 0, 0, 0, 0, 1, 1),
		(drawing, 2202, 2202, 0, 0, 0, 0, 1, 1),
		(drawing, 2201, 2201, 0, 0, 0, 0, 1, 1),
		(drawing, 2200, 2200, 0, 0, 0, 0, 1, 1),
		(drawing, 2199, 2199, 0, 0, 0, 0, 1, 1),
		(drawing, 2198, 2198, 0, 0, 0, 0, 1, 1),
		(drawing, 2197, 2197, 0, 0, 0, 0, 1, 1),
		(drawing, 2196, 2196, 0, 0, 0, 0, 1, 1),
		(drawing, 2195, 2195, 0, 0, 0, 0, 1, 1),
		(drawing, 2194, 2194, 0, 0, 0, 0, 1, 1),
		(drawing, 2193, 2193, 0, 0, 0, 0, 1, 1),
		(drawing, 2192, 2192, 0, 0, 0, 0, 1, 1),
		(drawing, 2191, 2191, 0, 0, 0, 0, 1, 1),
		(drawing, 2190, 2190, 0, 0, 0, 0, 1, 1),
		(drawing, 2189, 2189, 0, 0, 0, 0, 1, 1),
		(drawing, 2188, 2188, 0, 0, 0, 0, 1, 1),
		(drawing, 2187, 2187, 0, 0, 0, 0, 1, 1),
		(drawing, 2186, 2186, 0, 0, 0, 0, 1, 1),
		(drawing, 2185, 2185, 0, 0, 0, 0, 1, 1),
		(drawing, 2184, 2184, 0, 0, 0, 0, 1, 1),
		(drawing, 2183, 2183, 0, 0, 0, 0, 1, 1),
		(drawing, 2182, 2182, 0, 0, 0, 0, 1, 1),
		(drawing, 2181, 2181, 0, 0, 0, 0, 1, 1),
		(drawing, 2180, 2180, 0, 0, 0, 0, 1, 1),
		(drawing, 2179, 2179, 0, 0, 0, 0, 1, 1),
		(drawing, 2178, 2178, 0, 0, 0, 0, 1, 1),
		(drawing, 2177, 2177, 0, 0, 0, 0, 1, 1),
		(drawing, 2176, 2176, 0, 0, 0, 0, 1, 1),
		(drawing, 2175, 2175, 0, 0, 0, 0, 1, 1),
		(drawing, 2174, 2174, 0, 0, 0, 0, 1, 1),
		(drawing, 2173, 2173, 0, 0, 0, 0, 1, 1),
		(drawing, 2172, 2172, 0, 0, 0, 0, 1, 1),
		(drawing, 2171, 2171, 0, 0, 0, 0, 1, 1),
		(drawing, 2170, 2170, 0, 0, 0, 0, 1, 1),
		(drawing, 2169, 2169, 0, 0, 0, 0, 1, 1),
		(drawing, 2168, 2168, 0, 0, 0, 0, 1, 1),
		(drawing, 2167, 2167, 0, 0, 0, 0, 1, 1),
		(drawing, 2166, 2166, 0, 0, 0, 0, 1, 1),
		(drawing, 2165, 2165, 0, 0, 0, 0, 1, 1),
		(drawing, 2164, 2164, 0, 0, 0, 0, 1, 1),
		(drawing, 2163, 2163, 0, 0, 0, 0, 1, 1),
		(drawing, 2162, 2162, 0, 0, 0, 0, 1, 1),
		(drawing, 2161, 2161, 0, 0, 0, 0, 1, 1),
		(drawing, 2160, 2160, 0, 0, 0, 0, 1, 1),
		(drawing, 2159, 2159, 0, 0, 0, 0, 1, 1),
		(drawing, 2158, 2158, 0, 0, 0, 0, 1, 1),
		(drawing, 2157, 2157, 0, 0, 0, 0, 1, 1),
		(drawing, 2156, 2156, 0, 0, 0, 0, 1, 1),
		(drawing, 2155, 2155, 0, 0, 0, 0, 1, 1),
		(drawing, 2154, 2154, 0, 0, 0, 0, 1, 1),
		(drawing, 2153, 2153, 0, 0, 0, 0, 1, 1),
		(drawing, 2152, 2152, 0, 0, 0, 0, 1, 1),
		(drawing, 2151, 2151, 0, 0, 0, 0, 1, 1),
		(drawing, 2150, 2150, 0, 0, 0, 0, 1, 1),
		(drawing, 2149, 2149, 0, 0, 0, 0, 1, 1),
		(drawing, 2148, 2148, 0, 0, 0, 0, 1, 1),
		(drawing, 2147, 2147, 0, 0, 0, 0, 1, 1),
		(drawing, 2146, 2146, 0, 0, 0, 0, 1, 1),
		(drawing, 2145, 2145, 0, 0, 0, 0, 1, 1),
		(drawing, 2144, 2144, 0, 0, 0, 0, 1, 1),
		(drawing, 2143, 2143, 0, 0, 0, 0, 1, 1),
		(drawing, 2142, 2142, 0, 0, 0, 0, 1, 1),
		(drawing, 2141, 2141, 0, 0, 0, 0, 1, 1),
		(drawing, 2140, 2140, 0, 0, 0, 0, 1, 1),
		(drawing, 2139, 2139, 0, 0, 0, 0, 1, 1),
		(drawing, 2138, 2138, 0, 0, 0, 0, 1, 1),
		(drawing, 2137, 2137, 0, 0, 0, 0, 1, 1),
		(drawing, 2136, 2136, 0, 0, 0, 0, 1, 1),
		(drawing, 2135, 2135, 0, 0, 0, 0, 1, 1),
		(drawing, 2134, 2134, 0, 0, 0, 0, 1, 1),
		(drawing, 2133, 2133, 0, 0, 0, 0, 1, 1),
		(drawing, 2132, 2132, 0, 0, 0, 0, 1, 1),
		(drawing, 2131, 2131, 0, 0, 0, 0, 1, 1),
		(drawing, 2130, 2130, 0, 0, 0, 0, 1, 1),
		(drawing, 2129, 2129, 0, 0, 0, 0, 1, 1),
		(drawing, 2128, 2128, 0, 0, 0, 0, 1, 1),
		(drawing, 2127, 2127, 0, 0, 0, 0, 1, 1),
		(drawing, 2126, 2126, 0, 0, 0, 0, 1, 1),
		(drawing, 2125, 2125, 0, 0, 0, 0, 1, 1),
		(drawing, 2124, 2124, 0, 0, 0, 0, 1, 1),
		(drawing, 2123, 2123, 0, 0, 0, 0, 1, 1),
		(drawing, 2122, 2122, 0, 0, 0, 0, 1, 1),
		(drawing, 2121, 2121, 0, 0, 0, 0, 1, 1),
		(drawing, 2120, 2120, 0, 0, 0, 0, 1, 1),
		(drawing, 2119, 2119, 0, 0, 0, 0, 1, 1),
		(drawing, 2118, 2118, 0, 0, 0, 0, 1, 1),
		(drawing, 2117, 2117, 0, 0, 0, 0, 1, 1),
		(drawing, 2116, 2116, 0, 0, 0, 0, 1, 1),
		(drawing, 2115, 2115, 0, 0, 0, 0, 1, 1),
		(drawing, 2114, 2114, 0, 0, 0, 0, 1, 1),
		(drawing, 2113, 2113, 0, 0, 0, 0, 1, 1),
		(drawing, 2112, 2112, 0, 0, 0, 0, 1, 1),
		(drawing, 2111, 2111, 0, 0, 0, 0, 1, 1),
		(drawing, 2110, 2110, 0, 0, 0, 0, 1, 1),
		(drawing, 2109, 2109, 0, 0, 0, 0, 1, 1),
		(drawing, 2108, 2108, 0, 0, 0, 0, 1, 1),
		(drawing, 2107, 2107, 0, 0, 0, 0, 1, 1),
		(drawing, 2106, 2106, 0, 0, 0, 0, 1, 1),
		(drawing, 2105, 2105, 0, 0, 0, 0, 1, 1),
		(drawing, 2104, 2104, 0, 0, 0, 0, 1, 1),
		(drawing, 2103, 2103, 0, 0, 0, 0, 1, 1),
		(drawing, 2102, 2102, 0, 0, 0, 0, 1, 1),
		(drawing, 2101, 2101, 0, 0, 0, 0, 1, 1),
		(drawing, 2100, 2100, 0, 0, 0, 0, 1, 1),
		(drawing, 2099, 2099, 0, 0, 0, 0, 1, 1),
		(drawing, 2098, 2098, 0, 0, 0, 0, 1, 1),
		(drawing, 2097, 2097, 0, 0, 0, 0, 1, 1),
		(drawing, 2096, 2096, 0, 0, 0, 0, 1, 1),
		(drawing, 2095, 2095, 0, 0, 0, 0, 1, 1),
		(drawing, 2094, 2094, 0, 0, 0, 0, 1, 1),
		(drawing, 2093, 2093, 0, 0, 0, 0, 1, 1),
		(drawing, 2092, 2092, 0, 0, 0, 0, 1, 1),
		(drawing, 2091, 2091, 0, 0, 0, 0, 1, 1),
		(drawing, 2090, 2090, 0, 0, 0, 0, 1, 1),
		(drawing, 2089, 2089, 0, 0, 0, 0, 1, 1),
		(drawing, 2088, 2088, 0, 0, 0, 0, 1, 1),
		(drawing, 2087, 2087, 0, 0, 0, 0, 1, 1),
		(drawing, 2086, 2086, 0, 0, 0, 0, 1, 1),
		(drawing, 2085, 2085, 0, 0, 0, 0, 1, 1),
		(drawing, 2084, 2084, 0, 0, 0, 0, 1, 1),
		(drawing, 2083, 2083, 0, 0, 0, 0, 1, 1),
		(drawing, 2082, 2082, 0, 0, 0, 0, 1, 1),
		(drawing, 2081, 2081, 0, 0, 0, 0, 1, 1),
		(drawing, 2080, 2080, 0, 0, 0, 0, 1, 1),
		(drawing, 2079, 2079, 0, 0, 0, 0, 1, 1),
		(drawing, 2078, 2078, 0, 0, 0, 0, 1, 1),
		(drawing, 2077, 2077, 0, 0, 0, 0, 1, 1),
		(drawing, 2076, 2076, 0, 0, 0, 0, 1, 1),
		(drawing, 2075, 2075, 0, 0, 0, 0, 1, 1),
		(drawing, 2074, 2074, 0, 0, 0, 0, 1, 1),
		(drawing, 2073, 2073, 0, 0, 0, 0, 1, 1),
		(drawing, 2072, 2072, 0, 0, 0, 0, 1, 1),
		(drawing, 2071, 2071, 0, 0, 0, 0, 1, 1),
		(drawing, 2070, 2070, 0, 0, 0, 0, 1, 1),
		(drawing, 2069, 2069, 0, 0, 0, 0, 1, 1),
		(drawing, 2068, 2068, 0, 0, 0, 0, 1, 1),
		(drawing, 2067, 2067, 0, 0, 0, 0, 1, 1),
		(drawing, 2066, 2066, 0, 0, 0, 0, 1, 1),
		(drawing, 2065, 2065, 0, 0, 0, 0, 1, 1),
		(drawing, 2064, 2064, 0, 0, 0, 0, 1, 1),
		(drawing, 2063, 2063, 0, 0, 0, 0, 1, 1),
		(drawing, 2062, 2062, 0, 0, 0, 0, 1, 1),
		(drawing, 2061, 2061, 0, 0, 0, 0, 1, 1),
		(drawing, 2060, 2060, 0, 0, 0, 0, 1, 1),
		(drawing, 2059, 2059, 0, 0, 0, 0, 1, 1),
		(drawing, 2058, 2058, 0, 0, 0, 0, 1, 1),
		(drawing, 2057, 2057, 0, 0, 0, 0, 1, 1),
		(drawing, 2056, 2056, 0, 0, 0, 0, 1, 1),
		(drawing, 2055, 2055, 0, 0, 0, 0, 1, 1),
		(drawing, 2054, 2054, 0, 0, 0, 0, 1, 1),
		(drawing, 2053, 2053, 0, 0, 0, 0, 1, 1),
		(drawing, 2052, 2052, 0, 0, 0, 0, 1, 1),
		(drawing, 2051, 2051, 0, 0, 0, 0, 1, 1),
		(drawing, 2050, 2050, 0, 0, 0, 0, 1, 1),
		(drawing, 2049, 2049, 0, 0, 0, 0, 1, 1),
		(drawing, 2048, 2048, 0, 0, 0, 0, 1, 1),
		(drawing, 2047, 2047, 0, 0, 0, 0, 1, 1),
		(drawing, 2046, 2046, 0, 0, 0, 0, 1, 1),
		(drawing, 2045, 2045, 0, 0, 0, 0, 1, 1),
		(drawing, 2044, 2044, 0, 0, 0, 0, 1, 1),
		(drawing, 2043, 2043, 0, 0, 0, 0, 1, 1),
		(drawing, 2042, 2042, 0, 0, 0, 0, 1, 1),
		(drawing, 2041, 2041, 0, 0, 0, 0, 1, 1),
		(drawing, 2040, 2040, 0, 0, 0, 0, 1, 1),
		(drawing, 2039, 2039, 0, 0, 0, 0, 1, 1),
		(drawing, 2038, 2038, 0, 0, 0, 0, 1, 1),
		(drawing, 2037, 2037, 0, 0, 0, 0, 1, 1),
		(drawing, 2036, 2036, 0, 0, 0, 0, 1, 1),
		(drawing, 2035, 2035, 0, 0, 0, 0, 1, 1),
		(drawing, 2034, 2034, 0, 0, 0, 0, 1, 1),
		(drawing, 2033, 2033, 0, 0, 0, 0, 1, 1),
		(drawing, 2032, 2032, 0, 0, 0, 0, 1, 1),
		(drawing, 2031, 2031, 0, 0, 0, 0, 1, 1),
		(drawing, 2030, 2030, 0, 0, 0, 0, 1, 1),
		(drawing, 2029, 2029, 0, 0, 0, 0, 1, 1),
		(drawing, 2028, 2028, 0, 0, 0, 0, 1, 1),
		(drawing, 2027, 2027, 0, 0, 0, 0, 1, 1),
		(drawing, 2026, 2026, 0, 0, 0, 0, 1, 1),
		(drawing, 2025, 2025, 0, 0, 0, 0, 1, 1),
		(drawing, 2024, 2024, 0, 0, 0, 0, 1, 1),
		(drawing, 2023, 2023, 0, 0, 0, 0, 1, 1),
		(drawing, 2022, 2022, 0, 0, 0, 0, 1, 1),
		(drawing, 2021, 2021, 0, 0, 0, 0, 1, 1),
		(drawing, 2020, 2020, 0, 0, 0, 0, 1, 1),
		(drawing, 2019, 2019, 0, 0, 0, 0, 1, 1),
		(drawing, 2018, 2018, 0, 0, 0, 0, 1, 1),
		(drawing, 2017, 2017, 0, 0, 0, 0, 1, 1),
		(drawing, 2016, 2016, 0, 0, 0, 0, 1, 1),
		(drawing, 2015, 2015, 0, 0, 0, 0, 1, 1),
		(drawing, 2014, 2014, 0, 0, 0, 0, 1, 1),
		(drawing, 2013, 2013, 0, 0, 0, 0, 1, 1),
		(drawing, 2012, 2012, 0, 0, 0, 0, 1, 1),
		(drawing, 2011, 2011, 0, 0, 0, 0, 1, 1),
		(drawing, 2010, 2010, 0, 0, 0, 0, 1, 1),
		(drawing, 2009, 2009, 0, 0, 0, 0, 1, 1),
		(drawing, 2008, 2008, 0, 0, 0, 0, 1, 1),
		(drawing, 2007, 2007, 0, 0, 0, 0, 1, 1),
		(drawing, 2006, 2006, 0, 0, 0, 0, 1, 1),
		(drawing, 2005, 2005, 0, 0, 0, 0, 1, 1),
		(drawing, 2004, 2004, 0, 0, 0, 0, 1, 1),
		(drawing, 2003, 2003, 0, 0, 0, 0, 1, 1),
		(drawing, 2002, 2002, 0, 0, 0, 0, 1, 1),
		(drawing, 2001, 2001, 0, 0, 0, 0, 1, 1),
		(drawing, 2000, 2000, 0, 0, 0, 0, 1, 1),
		(drawing, 1999, 1999, 0, 0, 0, 0, 1, 1),
		(drawing, 1998, 1998, 0, 0, 0, 0, 1, 1),
		(drawing, 1997, 1997, 0, 0, 0, 0, 1, 1),
		(drawing, 1996, 1996, 0, 0, 0, 0, 1, 1),
		(drawing, 1995, 1995, 0, 0, 0, 0, 1, 1),
		(drawing, 1994, 1994, 0, 0, 0, 0, 1, 1),
		(drawing, 1993, 1993, 0, 0, 0, 0, 1, 1),
		(drawing, 1992, 1992, 0, 0, 0, 0, 1, 1),
		(drawing, 1991, 1991, 0, 0, 0, 0, 1, 1),
		(drawing, 1990, 1990, 0, 0, 0, 0, 1, 1),
		(drawing, 1989, 1989, 0, 0, 0, 0, 1, 1),
		(drawing, 1988, 1988, 0, 0, 0, 0, 1, 1),
		(drawing, 1987, 1987, 0, 0, 0, 0, 1, 1),
		(drawing, 1986, 1986, 0, 0, 0, 0, 1, 1),
		(drawing, 1985, 1985, 0, 0, 0, 0, 1, 1),
		(drawing, 1984, 1984, 0, 0, 0, 0, 1, 1),
		(drawing, 1983, 1983, 0, 0, 0, 0, 1, 1),
		(drawing, 1982, 1982, 0, 0, 0, 0, 1, 1),
		(drawing, 1981, 1981, 0, 0, 0, 0, 1, 1),
		(drawing, 1980, 1980, 0, 0, 0, 0, 1, 1),
		(drawing, 1979, 1979, 0, 0, 0, 0, 1, 1),
		(drawing, 1978, 1978, 0, 0, 0, 0, 1, 1),
		(drawing, 1977, 1977, 0, 0, 0, 0, 1, 1),
		(drawing, 1976, 1976, 0, 0, 0, 0, 1, 1),
		(drawing, 1975, 1975, 0, 0, 0, 0, 1, 1),
		(drawing, 1974, 1974, 0, 0, 0, 0, 1, 1),
		(drawing, 1973, 1973, 0, 0, 0, 0, 1, 1),
		(drawing, 1972, 1972, 0, 0, 0, 0, 1, 1),
		(drawing, 1971, 1971, 0, 0, 0, 0, 1, 1),
		(drawing, 1970, 1970, 0, 0, 0, 0, 1, 1),
		(drawing, 1969, 1969, 0, 0, 0, 0, 1, 1),
		(drawing, 1968, 1968, 0, 0, 0, 0, 1, 1),
		(drawing, 1967, 1967, 0, 0, 0, 0, 1, 1),
		(drawing, 1966, 1966, 0, 0, 0, 0, 1, 1),
		(drawing, 1965, 1965, 0, 0, 0, 0, 1, 1),
		(drawing, 1964, 1964, 0, 0, 0, 0, 1, 1),
		(drawing, 1963, 1963, 0, 0, 0, 0, 1, 1),
		(drawing, 1962, 1962, 0, 0, 0, 0, 1, 1),
		(drawing, 1961, 1961, 0, 0, 0, 0, 1, 1),
		(drawing, 1960, 1960, 0, 0, 0, 0, 1, 1),
		(drawing, 1959, 1959, 0, 0, 0, 0, 1, 1),
		(drawing, 1958, 1958, 0, 0, 0, 0, 1, 1),
		(drawing, 1957, 1957, 0, 0, 0, 0, 1, 1),
		(drawing, 1956, 1956, 0, 0, 0, 0, 1, 1),
		(drawing, 1955, 1955, 0, 0, 0, 0, 1, 1),
		(drawing, 1954, 1954, 0, 0, 0, 0, 1, 1),
		(drawing, 1953, 1953, 0, 0, 0, 0, 1, 1),
		(drawing, 1952, 1952, 0, 0, 0, 0, 1, 1),
		(drawing, 1951, 1951, 0, 0, 0, 0, 1, 1),
		(drawing, 1950, 1950, 0, 0, 0, 0, 1, 1),
		(drawing, 1949, 1949, 0, 0, 0, 0, 1, 1),
		(drawing, 1948, 1948, 0, 0, 0, 0, 1, 1),
		(drawing, 1947, 1947, 0, 0, 0, 0, 1, 1),
		(drawing, 1946, 1946, 0, 0, 0, 0, 1, 1),
		(drawing, 1945, 1945, 0, 0, 0, 0, 1, 1),
		(drawing, 1944, 1944, 0, 0, 0, 0, 1, 1),
		(drawing, 1943, 1943, 0, 0, 0, 0, 1, 1),
		(drawing, 1942, 1942, 0, 0, 0, 0, 1, 1),
		(drawing, 1941, 1941, 0, 0, 0, 0, 1, 1),
		(drawing, 1940, 1940, 0, 0, 0, 0, 1, 1),
		(drawing, 1939, 1939, 0, 0, 0, 0, 1, 1),
		(drawing, 1938, 1938, 0, 0, 0, 0, 1, 1),
		(drawing, 1937, 1937, 0, 0, 0, 0, 1, 1),
		(drawing, 1936, 1936, 0, 0, 0, 0, 1, 1),
		(drawing, 1935, 1935, 0, 0, 0, 0, 1, 1),
		(drawing, 1934, 1934, 0, 0, 0, 0, 1, 1),
		(drawing, 1933, 1933, 0, 0, 0, 0, 1, 1),
		(drawing, 1932, 1932, 0, 0, 0, 0, 1, 1),
		(drawing, 1931, 1931, 0, 0, 0, 0, 1, 1),
		(drawing, 1930, 1930, 0, 0, 0, 0, 1, 1),
		(drawing, 1929, 1929, 0, 0, 0, 0, 1, 1),
		(drawing, 1928, 1928, 0, 0, 0, 0, 1, 1),
		(drawing, 1927, 1927, 0, 0, 0, 0, 1, 1),
		(drawing, 1926, 1926, 0, 0, 0, 0, 1, 1),
		(drawing, 1925, 1925, 0, 0, 0, 0, 1, 1),
		(drawing, 1924, 1924, 0, 0, 0, 0, 1, 1),
		(drawing, 1923, 1923, 0, 0, 0, 0, 1, 1),
		(drawing, 1922, 1922, 0, 0, 0, 0, 1, 1),
		(drawing, 1921, 1921, 0, 0, 0, 0, 1, 1),
		(drawing, 1920, 1920, 0, 0, 0, 0, 1, 1),
		(drawing, 1919, 1919, 0, 0, 0, 0, 1, 1),
		(drawing, 1918, 1918, 0, 0, 0, 0, 1, 1),
		(drawing, 1917, 1917, 0, 0, 0, 0, 1, 1),
		(drawing, 1916, 1916, 0, 0, 0, 0, 1, 1),
		(drawing, 1915, 1915, 0, 0, 0, 0, 1, 1),
		(drawing, 1914, 1914, 0, 0, 0, 0, 1, 1),
		(drawing, 1913, 1913, 0, 0, 0, 0, 1, 1),
		(drawing, 1912, 1912, 0, 0, 0, 0, 1, 1),
		(drawing, 1911, 1911, 0, 0, 0, 0, 1, 1),
		(drawing, 1910, 1910, 0, 0, 0, 0, 1, 1),
		(drawing, 1909, 1909, 0, 0, 0, 0, 1, 1),
		(drawing, 1908, 1908, 0, 0, 0, 0, 1, 1),
		(drawing, 1907, 1907, 0, 0, 0, 0, 1, 1),
		(drawing, 1906, 1906, 0, 0, 0, 0, 1, 1),
		(drawing, 1905, 1905, 0, 0, 0, 0, 1, 1),
		(drawing, 1904, 1904, 0, 0, 0, 0, 1, 1),
		(drawing, 1903, 1903, 0, 0, 0, 0, 1, 1),
		(drawing, 1902, 1902, 0, 0, 0, 0, 1, 1),
		(drawing, 1901, 1901, 0, 0, 0, 0, 1, 1),
		(drawing, 1900, 1900, 0, 0, 0, 0, 1, 1),
		(drawing, 1899, 1899, 0, 0, 0, 0, 1, 1),
		(drawing, 1898, 1898, 0, 0, 0, 0, 1, 1),
		(drawing, 1897, 1897, 0, 0, 0, 0, 1, 1),
		(drawing, 1896, 1896, 0, 0, 0, 0, 1, 1),
		(drawing, 1895, 1895, 0, 0, 0, 0, 1, 1),
		(drawing, 1894, 1894, 0, 0, 0, 0, 1, 1),
		(drawing, 1893, 1893, 0, 0, 0, 0, 1, 1),
		(drawing, 1892, 1892, 0, 0, 0, 0, 1, 1),
		(drawing, 1891, 1891, 0, 0, 0, 0, 1, 1),
		(drawing, 1890, 1890, 0, 0, 0, 0, 1, 1),
		(drawing, 1889, 1889, 0, 0, 0, 0, 1, 1),
		(drawing, 1888, 1888, 0, 0, 0, 0, 1, 1),
		(drawing, 1887, 1887, 0, 0, 0, 0, 1, 1),
		(drawing, 1886, 1886, 0, 0, 0, 0, 1, 1),
		(drawing, 1885, 1885, 0, 0, 0, 0, 1, 1),
		(drawing, 1884, 1884, 0, 0, 0, 0, 1, 1),
		(drawing, 1883, 1883, 0, 0, 0, 0, 1, 1),
		(drawing, 1882, 1882, 0, 0, 0, 0, 1, 1),
		(drawing, 1881, 1881, 0, 0, 0, 0, 1, 1),
		(drawing, 1880, 1880, 0, 0, 0, 0, 1, 1),
		(drawing, 1879, 1879, 0, 0, 0, 0, 1, 1),
		(drawing, 1878, 1878, 0, 0, 0, 0, 1, 1),
		(drawing, 1877, 1877, 0, 0, 0, 0, 1, 1),
		(drawing, 1876, 1876, 0, 0, 0, 0, 1, 1),
		(drawing, 1875, 1875, 0, 0, 0, 0, 1, 1),
		(drawing, 1874, 1874, 0, 0, 0, 0, 1, 1),
		(drawing, 1873, 1873, 0, 0, 0, 0, 1, 1),
		(drawing, 1872, 1872, 0, 0, 0, 0, 1, 1),
		(drawing, 1871, 1871, 0, 0, 0, 0, 1, 1),
		(drawing, 1870, 1870, 0, 0, 0, 0, 1, 1),
		(drawing, 1869, 1869, 0, 0, 0, 0, 1, 1),
		(drawing, 1868, 1868, 0, 0, 0, 0, 1, 1),
		(drawing, 1867, 1867, 0, 0, 0, 0, 1, 1),
		(drawing, 1866, 1866, 0, 0, 0, 0, 1, 1),
		(drawing, 1865, 1865, 0, 0, 0, 0, 1, 1),
		(drawing, 1864, 1864, 0, 0, 0, 0, 1, 1),
		(drawing, 1863, 1863, 0, 0, 0, 0, 1, 1),
		(drawing, 1862, 1862, 0, 0, 0, 0, 1, 1),
		(drawing, 1861, 1861, 0, 0, 0, 0, 1, 1),
		(drawing, 1860, 1860, 0, 0, 0, 0, 1, 1),
		(drawing, 1859, 1859, 0, 0, 0, 0, 1, 1),
		(drawing, 1858, 1858, 0, 0, 0, 0, 1, 1),
		(drawing, 1857, 1857, 0, 0, 0, 0, 1, 1),
		(drawing, 1856, 1856, 0, 0, 0, 0, 1, 1),
		(drawing, 1855, 1855, 0, 0, 0, 0, 1, 1),
		(drawing, 1854, 1854, 0, 0, 0, 0, 1, 1),
		(drawing, 1853, 1853, 0, 0, 0, 0, 1, 1),
		(drawing, 1852, 1852, 0, 0, 0, 0, 1, 1),
		(drawing, 1851, 1851, 0, 0, 0, 0, 1, 1),
		(drawing, 1850, 1850, 0, 0, 0, 0, 1, 1),
		(drawing, 1849, 1849, 0, 0, 0, 0, 1, 1),
		(drawing, 1848, 1848, 0, 0, 0, 0, 1, 1),
		(drawing, 1847, 1847, 0, 0, 0, 0, 1, 1),
		(drawing, 1846, 1846, 0, 0, 0, 0, 1, 1),
		(drawing, 1845, 1845, 0, 0, 0, 0, 1, 1),
		(drawing, 1844, 1844, 0, 0, 0, 0, 1, 1),
		(drawing, 1843, 1843, 0, 0, 0, 0, 1, 1),
		(drawing, 1842, 1842, 0, 0, 0, 0, 1, 1),
		(drawing, 1841, 1841, 0, 0, 0, 0, 1, 1),
		(drawing, 1840, 1840, 0, 0, 0, 0, 1, 1),
		(drawing, 1839, 1839, 0, 0, 0, 0, 1, 1),
		(drawing, 1838, 1838, 0, 0, 0, 0, 1, 1),
		(drawing, 1837, 1837, 0, 0, 0, 0, 1, 1),
		(drawing, 1836, 1836, 0, 0, 0, 0, 1, 1),
		(drawing, 1835, 1835, 0, 0, 0, 0, 1, 1),
		(drawing, 1834, 1834, 0, 0, 0, 0, 1, 1),
		(drawing, 1833, 1833, 0, 0, 0, 0, 1, 1),
		(drawing, 1832, 1832, 0, 0, 0, 0, 1, 1),
		(drawing, 1831, 1831, 0, 0, 0, 0, 1, 1),
		(drawing, 1830, 1830, 0, 0, 0, 0, 1, 1),
		(drawing, 1829, 1829, 0, 0, 0, 0, 1, 1),
		(drawing, 1828, 1828, 0, 0, 0, 0, 1, 1),
		(drawing, 1827, 1827, 0, 0, 0, 0, 1, 1),
		(drawing, 1826, 1826, 0, 0, 0, 0, 1, 1),
		(drawing, 1825, 1825, 0, 0, 0, 0, 1, 1),
		(drawing, 1824, 1824, 0, 0, 0, 0, 1, 1),
		(drawing, 1823, 1823, 0, 0, 0, 0, 1, 1),
		(drawing, 1822, 1822, 0, 0, 0, 0, 1, 1),
		(drawing, 1821, 1821, 0, 0, 0, 0, 1, 1),
		(drawing, 1820, 1820, 0, 0, 0, 0, 1, 1),
		(drawing, 1819, 1819, 0, 0, 0, 0, 1, 1),
		(drawing, 1818, 1818, 0, 0, 0, 0, 1, 1),
		(drawing, 1817, 1817, 0, 0, 0, 0, 1, 1),
		(drawing, 1816, 1816, 0, 0, 0, 0, 1, 1),
		(drawing, 1815, 1815, 0, 0, 0, 0, 1, 1),
		(drawing, 1814, 1814, 0, 0, 0, 0, 1, 1),
		(drawing, 1813, 1813, 0, 0, 0, 0, 1, 1),
		(drawing, 1812, 1812, 0, 0, 0, 0, 1, 1),
		(drawing, 1811, 1811, 0, 0, 0, 0, 1, 1),
		(drawing, 1810, 1810, 0, 0, 0, 0, 1, 1),
		(drawing, 1809, 1809, 0, 0, 0, 0, 1, 1),
		(drawing, 1808, 1808, 0, 0, 0, 0, 1, 1),
		(drawing, 1807, 1807, 0, 0, 0, 0, 1, 1),
		(drawing, 1806, 1806, 0, 0, 0, 0, 1, 1),
		(drawing, 1805, 1805, 0, 0, 0, 0, 1, 1),
		(drawing, 1804, 1804, 0, 0, 0, 0, 1, 1),
		(drawing, 1803, 1803, 0, 0, 0, 0, 1, 1),
		(drawing, 1802, 1802, 0, 0, 0, 0, 1, 1),
		(drawing, 1801, 1801, 0, 0, 0, 0, 1, 1),
		(drawing, 1800, 1800, 0, 0, 0, 0, 1, 1),
		(drawing, 1799, 1799, 0, 0, 0, 0, 1, 1),
		(drawing, 1798, 1798, 0, 0, 0, 0, 1, 1),
		(drawing, 1797, 1797, 0, 0, 0, 0, 1, 1),
		(drawing, 1796, 1796, 0, 0, 0, 0, 1, 1),
		(drawing, 1795, 1795, 0, 0, 0, 0, 1, 1),
		(drawing, 1794, 1794, 0, 0, 0, 0, 1, 1),
		(drawing, 1793, 1793, 0, 0, 0, 0, 1, 1),
		(drawing, 1792, 1792, 0, 0, 0, 0, 1, 1),
		(drawing, 1791, 1791, 0, 0, 0, 0, 1, 1),
		(drawing, 1790, 1790, 0, 0, 0, 0, 1, 1),
		(drawing, 1789, 1789, 0, 0, 0, 0, 1, 1),
		(drawing, 1788, 1788, 0, 0, 0, 0, 1, 1),
		(drawing, 1787, 1787, 0, 0, 0, 0, 1, 1),
		(drawing, 1786, 1786, 0, 0, 0, 0, 1, 1),
		(drawing, 1785, 1785, 0, 0, 0, 0, 1, 1),
		(drawing, 1784, 1784, 0, 0, 0, 0, 1, 1),
		(drawing, 1783, 1783, 0, 0, 0, 0, 1, 1),
		(drawing, 1782, 1782, 0, 0, 0, 0, 1, 1),
		(drawing, 1781, 1781, 0, 0, 0, 0, 1, 1),
		(drawing, 1780, 1780, 0, 0, 0, 0, 1, 1),
		(drawing, 1779, 1779, 0, 0, 0, 0, 1, 1),
		(drawing, 1778, 1778, 0, 0, 0, 0, 1, 1),
		(drawing, 1777, 1777, 0, 0, 0, 0, 1, 1),
		(drawing, 1776, 1776, 0, 0, 0, 0, 1, 1),
		(drawing, 1775, 1775, 0, 0, 0, 0, 1, 1),
		(drawing, 1774, 1774, 0, 0, 0, 0, 1, 1),
		(drawing, 1773, 1773, 0, 0, 0, 0, 1, 1),
		(drawing, 1772, 1772, 0, 0, 0, 0, 1, 1),
		(drawing, 1771, 1771, 0, 0, 0, 0, 1, 1),
		(drawing, 1770, 1770, 0, 0, 0, 0, 1, 1),
		(drawing, 1769, 1769, 0, 0, 0, 0, 1, 1),
		(drawing, 1768, 1768, 0, 0, 0, 0, 1, 1),
		(drawing, 1767, 1767, 0, 0, 0, 0, 1, 1),
		(drawing, 1766, 1766, 0, 0, 0, 0, 1, 1),
		(drawing, 1765, 1765, 0, 0, 0, 0, 1, 1),
		(drawing, 1764, 1764, 0, 0, 0, 0, 1, 1),
		(drawing, 1763, 1763, 0, 0, 0, 0, 1, 1),
		(drawing, 1762, 1762, 0, 0, 0, 0, 1, 1),
		(drawing, 1761, 1761, 0, 0, 0, 0, 1, 1),
		(drawing, 1760, 1760, 0, 0, 0, 0, 1, 1),
		(drawing, 1759, 1759, 0, 0, 0, 0, 1, 1),
		(drawing, 1758, 1758, 0, 0, 0, 0, 1, 1),
		(drawing, 1757, 1757, 0, 0, 0, 0, 1, 1),
		(drawing, 1756, 1756, 0, 0, 0, 0, 1, 1),
		(drawing, 1755, 1755, 0, 0, 0, 0, 1, 1),
		(drawing, 1754, 1754, 0, 0, 0, 0, 1, 1),
		(drawing, 1753, 1753, 0, 0, 0, 0, 1, 1),
		(drawing, 1752, 1752, 0, 0, 0, 0, 1, 1),
		(drawing, 1751, 1751, 0, 0, 0, 0, 1, 1),
		(drawing, 1750, 1750, 0, 0, 0, 0, 1, 1),
		(drawing, 1749, 1749, 0, 0, 0, 0, 1, 1),
		(drawing, 1748, 1748, 0, 0, 0, 0, 1, 1),
		(drawing, 1747, 1747, 0, 0, 0, 0, 1, 1),
		(drawing, 1746, 1746, 0, 0, 0, 0, 1, 1),
		(drawing, 1745, 1745, 0, 0, 0, 0, 1, 1),
		(drawing, 1744, 1744, 0, 0, 0, 0, 1, 1),
		(drawing, 1743, 1743, 0, 0, 0, 0, 1, 1),
		(drawing, 1742, 1742, 0, 0, 0, 0, 1, 1),
		(drawing, 1741, 1741, 0, 0, 0, 0, 1, 1),
		(drawing, 1740, 1740, 0, 0, 0, 0, 1, 1),
		(drawing, 1739, 1739, 0, 0, 0, 0, 1, 1),
		(drawing, 1738, 1738, 0, 0, 0, 0, 1, 1),
		(drawing, 1737, 1737, 0, 0, 0, 0, 1, 1),
		(drawing, 1736, 1736, 0, 0, 0, 0, 1, 1),
		(drawing, 1735, 1735, 0, 0, 0, 0, 1, 1),
		(drawing, 1734, 1734, 0, 0, 0, 0, 1, 1),
		(drawing, 1733, 1733, 0, 0, 0, 0, 1, 1),
		(drawing, 1732, 1732, 0, 0, 0, 0, 1, 1),
		(drawing, 1731, 1731, 0, 0, 0, 0, 1, 1),
		(drawing, 1730, 1730, 0, 0, 0, 0, 1, 1),
		(drawing, 1729, 1729, 0, 0, 0, 0, 1, 1),
		(drawing, 1728, 1728, 0, 0, 0, 0, 1, 1),
		(drawing, 1727, 1727, 0, 0, 0, 0, 1, 1),
		(drawing, 1726, 1726, 0, 0, 0, 0, 1, 1),
		(drawing, 1725, 1725, 0, 0, 0, 0, 1, 1),
		(drawing, 1724, 1724, 0, 0, 0, 0, 1, 1),
		(drawing, 1723, 1723, 0, 0, 0, 0, 1, 1),
		(drawing, 1722, 1722, 0, 0, 0, 0, 1, 1),
		(drawing, 1721, 1721, 0, 0, 0, 0, 1, 1),
		(drawing, 1720, 1720, 0, 0, 0, 0, 1, 1),
		(drawing, 1719, 1719, 0, 0, 0, 0, 1, 1),
		(drawing, 1718, 1718, 0, 0, 0, 0, 1, 1),
		(drawing, 1717, 1717, 0, 0, 0, 0, 1, 1),
		(drawing, 1716, 1716, 0, 0, 0, 0, 1, 1),
		(drawing, 1715, 1715, 0, 0, 0, 0, 1, 1),
		(drawing, 1714, 1714, 0, 0, 0, 0, 1, 1),
		(drawing, 1713, 1713, 0, 0, 0, 0, 1, 1),
		(drawing, 1712, 1712, 0, 0, 0, 0, 1, 1),
		(drawing, 1711, 1711, 0, 0, 0, 0, 1, 1),
		(drawing, 1710, 1710, 0, 0, 0, 0, 1, 1),
		(drawing, 1709, 1709, 0, 0, 0, 0, 1, 1),
		(drawing, 1708, 1708, 0, 0, 0, 0, 1, 1),
		(drawing, 1707, 1707, 0, 0, 0, 0, 1, 1),
		(drawing, 1706, 1706, 0, 0, 0, 0, 1, 1),
		(drawing, 1705, 1705, 0, 0, 0, 0, 1, 1),
		(drawing, 1704, 1704, 0, 0, 0, 0, 1, 1),
		(drawing, 1703, 1703, 0, 0, 0, 0, 1, 1),
		(drawing, 1702, 1702, 0, 0, 0, 0, 1, 1),
		(drawing, 1701, 1701, 0, 0, 0, 0, 1, 1),
		(drawing, 1700, 1700, 0, 0, 0, 0, 1, 1),
		(drawing, 1699, 1699, 0, 0, 0, 0, 1, 1),
		(drawing, 1698, 1698, 0, 0, 0, 0, 1, 1),
		(drawing, 1697, 1697, 0, 0, 0, 0, 1, 1),
		(drawing, 1696, 1696, 0, 0, 0, 0, 1, 1),
		(drawing, 1695, 1695, 0, 0, 0, 0, 1, 1),
		(drawing, 1694, 1694, 0, 0, 0, 0, 1, 1),
		(drawing, 1693, 1693, 0, 0, 0, 0, 1, 1),
		(drawing, 1692, 1692, 0, 0, 0, 0, 1, 1),
		(drawing, 1691, 1691, 0, 0, 0, 0, 1, 1),
		(drawing, 1690, 1690, 0, 0, 0, 0, 1, 1),
		(drawing, 1689, 1689, 0, 0, 0, 0, 1, 1),
		(drawing, 1688, 1688, 0, 0, 0, 0, 1, 1),
		(drawing, 1687, 1687, 0, 0, 0, 0, 1, 1),
		(drawing, 1686, 1686, 0, 0, 0, 0, 1, 1),
		(drawing, 1685, 1685, 0, 0, 0, 0, 1, 1),
		(drawing, 1684, 1684, 0, 0, 0, 0, 1, 1),
		(drawing, 1683, 1683, 0, 0, 0, 0, 1, 1),
		(drawing, 1682, 1682, 0, 0, 0, 0, 1, 1),
		(drawing, 1681, 1681, 0, 0, 0, 0, 1, 1),
		(drawing, 1680, 1680, 0, 0, 0, 0, 1, 1),
		(drawing, 1679, 1679, 0, 0, 0, 0, 1, 1),
		(drawing, 1678, 1678, 0, 0, 0, 0, 1, 1),
		(drawing, 1677, 1677, 0, 0, 0, 0, 1, 1),
		(drawing, 1676, 1676, 0, 0, 0, 0, 1, 1),
		(drawing, 1675, 1675, 0, 0, 0, 0, 1, 1),
		(drawing, 1674, 1674, 0, 0, 0, 0, 1, 1),
		(drawing, 1673, 1673, 0, 0, 0, 0, 1, 1),
		(drawing, 1672, 1672, 0, 0, 0, 0, 1, 1),
		(drawing, 1671, 1671, 0, 0, 0, 0, 1, 1),
		(drawing, 1670, 1670, 0, 0, 0, 0, 1, 1),
		(drawing, 1669, 1669, 0, 0, 0, 0, 1, 1),
		(drawing, 1668, 1668, 0, 0, 0, 0, 1, 1),
		(drawing, 1667, 1667, 0, 0, 0, 0, 1, 1),
		(drawing, 1666, 1666, 0, 0, 0, 0, 1, 1),
		(drawing, 1665, 1665, 0, 0, 0, 0, 1, 1),
		(drawing, 1664, 1664, 0, 0, 0, 0, 1, 1),
		(drawing, 1663, 1663, 0, 0, 0, 0, 1, 1),
		(drawing, 1662, 1662, 0, 0, 0, 0, 1, 1),
		(drawing, 1661, 1661, 0, 0, 0, 0, 1, 1),
		(drawing, 1660, 1660, 0, 0, 0, 0, 1, 1),
		(drawing, 1659, 1659, 0, 0, 0, 0, 1, 1),
		(drawing, 1658, 1658, 0, 0, 0, 0, 1, 1),
		(drawing, 1657, 1657, 0, 0, 0, 0, 1, 1),
		(drawing, 1656, 1656, 0, 0, 0, 0, 1, 1),
		(drawing, 1655, 1655, 0, 0, 0, 0, 1, 1),
		(drawing, 1654, 1654, 0, 0, 0, 0, 1, 1),
		(drawing, 1653, 1653, 0, 0, 0, 0, 1, 1),
		(drawing, 1652, 1652, 0, 0, 0, 0, 1, 1),
		(drawing, 1651, 1651, 0, 0, 0, 0, 1, 1),
		(drawing, 1650, 1650, 0, 0, 0, 0, 1, 1),
		(drawing, 1649, 1649, 0, 0, 0, 0, 1, 1),
		(drawing, 1648, 1648, 0, 0, 0, 0, 1, 1),
		(drawing, 1647, 1647, 0, 0, 0, 0, 1, 1),
		(drawing, 1646, 1646, 0, 0, 0, 0, 1, 1),
		(drawing, 1645, 1645, 0, 0, 0, 0, 1, 1),
		(drawing, 1644, 1644, 0, 0, 0, 0, 1, 1),
		(drawing, 1643, 1643, 0, 0, 0, 0, 1, 1),
		(drawing, 1642, 1642, 0, 0, 0, 0, 1, 1),
		(drawing, 1641, 1641, 0, 0, 0, 0, 1, 1),
		(drawing, 1640, 1640, 0, 0, 0, 0, 1, 1),
		(drawing, 1639, 1639, 0, 0, 0, 0, 1, 1),
		(drawing, 1638, 1638, 0, 0, 0, 0, 1, 1),
		(drawing, 1637, 1637, 0, 0, 0, 0, 1, 1),
		(drawing, 1636, 1636, 0, 0, 0, 0, 1, 1),
		(drawing, 1635, 1635, 0, 0, 0, 0, 1, 1),
		(drawing, 1634, 1634, 0, 0, 0, 0, 1, 1),
		(drawing, 1633, 1633, 0, 0, 0, 0, 1, 1),
		(drawing, 1632, 1632, 0, 0, 0, 0, 1, 1),
		(drawing, 1631, 1631, 0, 0, 0, 0, 1, 1),
		(drawing, 1630, 1630, 0, 0, 0, 0, 1, 1),
		(drawing, 1629, 1629, 0, 0, 0, 0, 1, 1),
		(drawing, 1628, 1628, 0, 0, 0, 0, 1, 1),
		(drawing, 1627, 1627, 0, 0, 0, 0, 1, 1),
		(drawing, 1626, 1626, 0, 0, 0, 0, 1, 1),
		(drawing, 1625, 1625, 0, 0, 0, 0, 1, 1),
		(drawing, 1624, 1624, 0, 0, 0, 0, 1, 1),
		(drawing, 1623, 1623, 0, 0, 0, 0, 1, 1),
		(drawing, 1622, 1622, 0, 0, 0, 0, 1, 1),
		(drawing, 1621, 1621, 0, 0, 0, 0, 1, 1),
		(drawing, 1620, 1620, 0, 0, 0, 0, 1, 1),
		(drawing, 1619, 1619, 0, 0, 0, 0, 1, 1),
		(drawing, 1618, 1618, 0, 0, 0, 0, 1, 1),
		(drawing, 1617, 1617, 0, 0, 0, 0, 1, 1),
		(drawing, 1616, 1616, 0, 0, 0, 0, 1, 1),
		(drawing, 1615, 1615, 0, 0, 0, 0, 1, 1),
		(drawing, 1614, 1614, 0, 0, 0, 0, 1, 1),
		(drawing, 1613, 1613, 0, 0, 0, 0, 1, 1),
		(drawing, 1612, 1612, 0, 0, 0, 0, 1, 1),
		(drawing, 1611, 1611, 0, 0, 0, 0, 1, 1),
		(drawing, 1610, 1610, 0, 0, 0, 0, 1, 1),
		(drawing, 1609, 1609, 0, 0, 0, 0, 1, 1),
		(drawing, 1608, 1608, 0, 0, 0, 0, 1, 1),
		(drawing, 1607, 1607, 0, 0, 0, 0, 1, 1),
		(drawing, 1606, 1606, 0, 0, 0, 0, 1, 1),
		(drawing, 1605, 1605, 0, 0, 0, 0, 1, 1),
		(drawing, 1604, 1604, 0, 0, 0, 0, 1, 1),
		(drawing, 1603, 1603, 0, 0, 0, 0, 1, 1),
		(drawing, 1602, 1602, 0, 0, 0, 0, 1, 1),
		(drawing, 1601, 1601, 0, 0, 0, 0, 1, 1),
		(drawing, 1600, 1600, 0, 0, 0, 0, 1, 1),
		(drawing, 1599, 1599, 0, 0, 0, 0, 1, 1),
		(drawing, 1598, 1598, 0, 0, 0, 0, 1, 1),
		(drawing, 1597, 1597, 0, 0, 0, 0, 1, 1),
		(drawing, 1596, 1596, 0, 0, 0, 0, 1, 1),
		(drawing, 1595, 1595, 0, 0, 0, 0, 1, 1),
		(drawing, 1594, 1594, 0, 0, 0, 0, 1, 1),
		(drawing, 1593, 1593, 0, 0, 0, 0, 1, 1),
		(drawing, 1592, 1592, 0, 0, 0, 0, 1, 1),
		(drawing, 1591, 1591, 0, 0, 0, 0, 1, 1),
		(drawing, 1590, 1590, 0, 0, 0, 0, 1, 1),
		(drawing, 1589, 1589, 0, 0, 0, 0, 1, 1),
		(drawing, 1588, 1588, 0, 0, 0, 0, 1, 1),
		(drawing, 1587, 1587, 0, 0, 0, 0, 1, 1),
		(drawing, 1586, 1586, 0, 0, 0, 0, 1, 1),
		(drawing, 1585, 1585, 0, 0, 0, 0, 1, 1),
		(drawing, 1584, 1584, 0, 0, 0, 0, 1, 1),
		(drawing, 1583, 1583, 0, 0, 0, 0, 1, 1),
		(drawing, 1582, 1582, 0, 0, 0, 0, 1, 1),
		(drawing, 1581, 1581, 0, 0, 0, 0, 1, 1),
		(drawing, 1580, 1580, 0, 0, 0, 0, 1, 1),
		(drawing, 1579, 1579, 0, 0, 0, 0, 1, 1),
		(drawing, 1578, 1578, 0, 0, 0, 0, 1, 1),
		(drawing, 1577, 1577, 0, 0, 0, 0, 1, 1),
		(drawing, 1576, 1576, 0, 0, 0, 0, 1, 1),
		(drawing, 1575, 1575, 0, 0, 0, 0, 1, 1),
		(drawing, 1574, 1574, 0, 0, 0, 0, 1, 1),
		(drawing, 1573, 1573, 0, 0, 0, 0, 1, 1),
		(drawing, 1572, 1572, 0, 0, 0, 0, 1, 1),
		(drawing, 1571, 1571, 0, 0, 0, 0, 1, 1),
		(drawing, 1570, 1570, 0, 0, 0, 0, 1, 1),
		(drawing, 1569, 1569, 0, 0, 0, 0, 1, 1),
		(drawing, 1568, 1568, 0, 0, 0, 0, 1, 1),
		(drawing, 1567, 1567, 0, 0, 0, 0, 1, 1),
		(drawing, 1566, 1566, 0, 0, 0, 0, 1, 1),
		(drawing, 1565, 1565, 0, 0, 0, 0, 1, 1),
		(drawing, 1564, 1564, 0, 0, 0, 0, 1, 1),
		(drawing, 1563, 1563, 0, 0, 0, 0, 1, 1),
		(drawing, 1562, 1562, 0, 0, 0, 0, 1, 1),
		(drawing, 1561, 1561, 0, 0, 0, 0, 1, 1),
		(drawing, 1560, 1560, 0, 0, 0, 0, 1, 1),
		(drawing, 1559, 1559, 0, 0, 0, 0, 1, 1),
		(drawing, 1558, 1558, 0, 0, 0, 0, 1, 1),
		(drawing, 1557, 1557, 0, 0, 0, 0, 1, 1),
		(drawing, 1556, 1556, 0, 0, 0, 0, 1, 1),
		(drawing, 1555, 1555, 0, 0, 0, 0, 1, 1),
		(drawing, 1554, 1554, 0, 0, 0, 0, 1, 1),
		(drawing, 1553, 1553, 0, 0, 0, 0, 1, 1),
		(drawing, 1552, 1552, 0, 0, 0, 0, 1, 1),
		(drawing, 1551, 1551, 0, 0, 0, 0, 1, 1),
		(drawing, 1550, 1550, 0, 0, 0, 0, 1, 1),
		(drawing, 1549, 1549, 0, 0, 0, 0, 1, 1),
		(drawing, 1548, 1548, 0, 0, 0, 0, 1, 1),
		(drawing, 1547, 1547, 0, 0, 0, 0, 1, 1),
		(drawing, 1546, 1546, 0, 0, 0, 0, 1, 1),
		(drawing, 1545, 1545, 0, 0, 0, 0, 1, 1),
		(drawing, 1544, 1544, 0, 0, 0, 0, 1, 1),
		(drawing, 1543, 1543, 0, 0, 0, 0, 1, 1),
		(drawing, 1542, 1542, 0, 0, 0, 0, 1, 1),
		(drawing, 1541, 1541, 0, 0, 0, 0, 1, 1),
		(drawing, 1540, 1540, 0, 0, 0, 0, 1, 1),
		(drawing, 1539, 1539, 0, 0, 0, 0, 1, 1),
		(drawing, 1538, 1538, 0, 0, 0, 0, 1, 1),
		(drawing, 1537, 1537, 0, 0, 0, 0, 1, 1),
		(drawing, 1536, 1536, 0, 0, 0, 0, 1, 1),
		(drawing, 1535, 1535, 0, 0, 0, 0, 1, 1),
		(drawing, 1534, 1534, 0, 0, 0, 0, 1, 1),
		(drawing, 1533, 1533, 0, 0, 0, 0, 1, 1),
		(drawing, 1532, 1532, 0, 0, 0, 0, 1, 1),
		(drawing, 1531, 1531, 0, 0, 0, 0, 1, 1),
		(drawing, 1530, 1530, 0, 0, 0, 0, 1, 1),
		(drawing, 1529, 1529, 0, 0, 0, 0, 1, 1),
		(drawing, 1528, 1528, 0, 0, 0, 0, 1, 1),
		(drawing, 1527, 1527, 0, 0, 0, 0, 1, 1),
		(drawing, 1526, 1526, 0, 0, 0, 0, 1, 1),
		(drawing, 1525, 1525, 0, 0, 0, 0, 1, 1),
		(drawing, 1524, 1524, 0, 0, 0, 0, 1, 1),
		(drawing, 1523, 1523, 0, 0, 0, 0, 1, 1),
		(drawing, 1522, 1522, 0, 0, 0, 0, 1, 1),
		(drawing, 1521, 1521, 0, 0, 0, 0, 1, 1),
		(drawing, 1520, 1520, 0, 0, 0, 0, 1, 1),
		(drawing, 1519, 1519, 0, 0, 0, 0, 1, 1),
		(drawing, 1518, 1518, 0, 0, 0, 0, 1, 1),
		(drawing, 1517, 1517, 0, 0, 0, 0, 1, 1),
		(drawing, 1516, 1516, 0, 0, 0, 0, 1, 1),
		(drawing, 1515, 1515, 0, 0, 0, 0, 1, 1),
		(drawing, 1514, 1514, 0, 0, 0, 0, 1, 1),
		(drawing, 1513, 1513, 0, 0, 0, 0, 1, 1),
		(drawing, 1512, 1512, 0, 0, 0, 0, 1, 1),
		(drawing, 1511, 1511, 0, 0, 0, 0, 1, 1),
		(drawing, 1510, 1510, 0, 0, 0, 0, 1, 1),
		(drawing, 1509, 1509, 0, 0, 0, 0, 1, 1),
		(drawing, 1508, 1508, 0, 0, 0, 0, 1, 1),
		(drawing, 1507, 1507, 0, 0, 0, 0, 1, 1),
		(drawing, 1506, 1506, 0, 0, 0, 0, 1, 1),
		(drawing, 1505, 1505, 0, 0, 0, 0, 1, 1),
		(drawing, 1504, 1504, 0, 0, 0, 0, 1, 1),
		(drawing, 1503, 1503, 0, 0, 0, 0, 1, 1),
		(drawing, 1502, 1502, 0, 0, 0, 0, 1, 1),
		(drawing, 1501, 1501, 0, 0, 0, 0, 1, 1),
		(drawing, 1500, 1500, 0, 0, 0, 0, 1, 1),
		(drawing, 1499, 1499, 0, 0, 0, 0, 1, 1),
		(drawing, 1498, 1498, 0, 0, 0, 0, 1, 1),
		(drawing, 1497, 1497, 0, 0, 0, 0, 1, 1),
		(drawing, 1496, 1496, 0, 0, 0, 0, 1, 1),
		(drawing, 1495, 1495, 0, 0, 0, 0, 1, 1),
		(drawing, 1494, 1494, 0, 0, 0, 0, 1, 1),
		(drawing, 1493, 1493, 0, 0, 0, 0, 1, 1),
		(drawing, 1492, 1492, 0, 0, 0, 0, 1, 1),
		(drawing, 1491, 1491, 0, 0, 0, 0, 1, 1),
		(drawing, 1490, 1490, 0, 0, 0, 0, 1, 1),
		(drawing, 1489, 1489, 0, 0, 0, 0, 1, 1),
		(drawing, 1488, 1488, 0, 0, 0, 0, 1, 1),
		(drawing, 1487, 1487, 0, 0, 0, 0, 1, 1),
		(drawing, 1486, 1486, 0, 0, 0, 0, 1, 1),
		(drawing, 1485, 1485, 0, 0, 0, 0, 1, 1),
		(drawing, 1484, 1484, 0, 0, 0, 0, 1, 1),
		(drawing, 1483, 1483, 0, 0, 0, 0, 1, 1),
		(drawing, 1482, 1482, 0, 0, 0, 0, 1, 1),
		(drawing, 1481, 1481, 0, 0, 0, 0, 1, 1),
		(drawing, 1480, 1480, 0, 0, 0, 0, 1, 1),
		(drawing, 1479, 1479, 0, 0, 0, 0, 1, 1),
		(drawing, 1478, 1478, 0, 0, 0, 0, 1, 1),
		(drawing, 1477, 1477, 0, 0, 0, 0, 1, 1),
		(drawing, 1476, 1476, 0, 0, 0, 0, 1, 1),
		(drawing, 1475, 1475, 0, 0, 0, 0, 1, 1),
		(drawing, 1474, 1474, 0, 0, 0, 0, 1, 1),
		(drawing, 1473, 1473, 0, 0, 0, 0, 1, 1),
		(drawing, 1472, 1472, 0, 0, 0, 0, 1, 1),
		(drawing, 1471, 1471, 0, 0, 0, 0, 1, 1),
		(drawing, 1470, 1470, 0, 0, 0, 0, 1, 1),
		(drawing, 1469, 1469, 0, 0, 0, 0, 1, 1),
		(drawing, 1468, 1468, 0, 0, 0, 0, 1, 1),
		(drawing, 1467, 1467, 0, 0, 0, 0, 1, 1),
		(drawing, 1466, 1466, 0, 0, 0, 0, 1, 1),
		(drawing, 1465, 1465, 0, 0, 0, 0, 1, 1),
		(drawing, 1464, 1464, 0, 0, 0, 0, 1, 1),
		(drawing, 1463, 1463, 0, 0, 0, 0, 1, 1),
		(drawing, 1462, 1462, 0, 0, 0, 0, 1, 1),
		(drawing, 1461, 1461, 0, 0, 0, 0, 1, 1),
		(drawing, 1460, 1460, 0, 0, 0, 0, 1, 1),
		(drawing, 1459, 1459, 0, 0, 0, 0, 1, 1),
		(drawing, 1458, 1458, 0, 0, 0, 0, 1, 1),
		(drawing, 1457, 1457, 0, 0, 0, 0, 1, 1),
		(drawing, 1456, 1456, 0, 0, 0, 0, 1, 1),
		(drawing, 1455, 1455, 0, 0, 0, 0, 1, 1),
		(drawing, 1454, 1454, 0, 0, 0, 0, 1, 1),
		(drawing, 1453, 1453, 0, 0, 0, 0, 1, 1),
		(drawing, 1452, 1452, 0, 0, 0, 0, 1, 1),
		(drawing, 1451, 1451, 0, 0, 0, 0, 1, 1),
		(drawing, 1450, 1450, 0, 0, 0, 0, 1, 1),
		(drawing, 1449, 1449, 0, 0, 0, 0, 1, 1),
		(drawing, 1448, 1448, 0, 0, 0, 0, 1, 1),
		(drawing, 1447, 1447, 0, 0, 0, 0, 1, 1),
		(drawing, 1446, 1446, 0, 0, 0, 0, 1, 1),
		(drawing, 1445, 1445, 0, 0, 0, 0, 1, 1),
		(drawing, 1444, 1444, 0, 0, 0, 0, 1, 1),
		(drawing, 1443, 1443, 0, 0, 0, 0, 1, 1),
		(drawing, 1442, 1442, 0, 0, 0, 0, 1, 1),
		(drawing, 1441, 1441, 0, 0, 0, 0, 1, 1),
		(drawing, 1440, 1440, 0, 0, 0, 0, 1, 1),
		(drawing, 1439, 1439, 0, 0, 0, 0, 1, 1),
		(drawing, 1438, 1438, 0, 0, 0, 0, 1, 1),
		(drawing, 1437, 1437, 0, 0, 0, 0, 1, 1),
		(drawing, 1436, 1436, 0, 0, 0, 0, 1, 1),
		(drawing, 1435, 1435, 0, 0, 0, 0, 1, 1),
		(drawing, 1434, 1434, 0, 0, 0, 0, 1, 1),
		(drawing, 1433, 1433, 0, 0, 0, 0, 1, 1),
		(drawing, 1432, 1432, 0, 0, 0, 0, 1, 1),
		(drawing, 1431, 1431, 0, 0, 0, 0, 1, 1),
		(drawing, 1430, 1430, 0, 0, 0, 0, 1, 1),
		(drawing, 1429, 1429, 0, 0, 0, 0, 1, 1),
		(drawing, 1428, 1428, 0, 0, 0, 0, 1, 1),
		(drawing, 1427, 1427, 0, 0, 0, 0, 1, 1),
		(drawing, 1426, 1426, 0, 0, 0, 0, 1, 1),
		(drawing, 1425, 1425, 0, 0, 0, 0, 1, 1),
		(drawing, 1424, 1424, 0, 0, 0, 0, 1, 1),
		(drawing, 1423, 1423, 0, 0, 0, 0, 1, 1),
		(drawing, 1422, 1422, 0, 0, 0, 0, 1, 1),
		(drawing, 1421, 1421, 0, 0, 0, 0, 1, 1),
		(drawing, 1420, 1420, 0, 0, 0, 0, 1, 1),
		(drawing, 1419, 1419, 0, 0, 0, 0, 1, 1),
		(drawing, 1418, 1418, 0, 0, 0, 0, 1, 1),
		(drawing, 1417, 1417, 0, 0, 0, 0, 1, 1),
		(drawing, 1416, 1416, 0, 0, 0, 0, 1, 1),
		(drawing, 1415, 1415, 0, 0, 0, 0, 1, 1),
		(drawing, 1414, 1414, 0, 0, 0, 0, 1, 1),
		(drawing, 1413, 1413, 0, 0, 0, 0, 1, 1),
		(drawing, 1412, 1412, 0, 0, 0, 0, 1, 1),
		(drawing, 1411, 1411, 0, 0, 0, 0, 1, 1),
		(drawing, 1410, 1410, 0, 0, 0, 0, 1, 1),
		(drawing, 1409, 1409, 0, 0, 0, 0, 1, 1),
		(drawing, 1408, 1408, 0, 0, 0, 0, 1, 1),
		(drawing, 1407, 1407, 0, 0, 0, 0, 1, 1),
		(drawing, 1406, 1406, 0, 0, 0, 0, 1, 1),
		(drawing, 1405, 1405, 0, 0, 0, 0, 1, 1),
		(drawing, 1404, 1404, 0, 0, 0, 0, 1, 1),
		(drawing, 1403, 1403, 0, 0, 0, 0, 1, 1),
		(drawing, 1402, 1402, 0, 0, 0, 0, 1, 1),
		(drawing, 1401, 1401, 0, 0, 0, 0, 1, 1),
		(drawing, 1400, 1400, 0, 0, 0, 0, 1, 1),
		(drawing, 1399, 1399, 0, 0, 0, 0, 1, 1),
		(drawing, 1398, 1398, 0, 0, 0, 0, 1, 1),
		(drawing, 1397, 1397, 0, 0, 0, 0, 1, 1),
		(drawing, 1396, 1396, 0, 0, 0, 0, 1, 1),
		(drawing, 1395, 1395, 0, 0, 0, 0, 1, 1),
		(drawing, 1394, 1394, 0, 0, 0, 0, 1, 1),
		(drawing, 1393, 1393, 0, 0, 0, 0, 1, 1),
		(drawing, 1392, 1392, 0, 0, 0, 0, 1, 1),
		(drawing, 1391, 1391, 0, 0, 0, 0, 1, 1),
		(drawing, 1390, 1390, 0, 0, 0, 0, 1, 1),
		(drawing, 1389, 1389, 0, 0, 0, 0, 1, 1),
		(drawing, 1388, 1388, 0, 0, 0, 0, 1, 1),
		(drawing, 1387, 1387, 0, 0, 0, 0, 1, 1),
		(drawing, 1386, 1386, 0, 0, 0, 0, 1, 1),
		(drawing, 1385, 1385, 0, 0, 0, 0, 1, 1),
		(drawing, 1384, 1384, 0, 0, 0, 0, 1, 1),
		(drawing, 1383, 1383, 0, 0, 0, 0, 1, 1),
		(drawing, 1382, 1382, 0, 0, 0, 0, 1, 1),
		(drawing, 1381, 1381, 0, 0, 0, 0, 1, 1),
		(drawing, 1380, 1380, 0, 0, 0, 0, 1, 1),
		(drawing, 1379, 1379, 0, 0, 0, 0, 1, 1),
		(drawing, 1378, 1378, 0, 0, 0, 0, 1, 1),
		(drawing, 1377, 1377, 0, 0, 0, 0, 1, 1),
		(drawing, 1376, 1376, 0, 0, 0, 0, 1, 1),
		(drawing, 1375, 1375, 0, 0, 0, 0, 1, 1),
		(drawing, 1374, 1374, 0, 0, 0, 0, 1, 1),
		(drawing, 1373, 1373, 0, 0, 0, 0, 1, 1),
		(drawing, 1372, 1372, 0, 0, 0, 0, 1, 1),
		(drawing, 1371, 1371, 0, 0, 0, 0, 1, 1),
		(drawing, 1370, 1370, 0, 0, 0, 0, 1, 1),
		(drawing, 1369, 1369, 0, 0, 0, 0, 1, 1),
		(drawing, 1368, 1368, 0, 0, 0, 0, 1, 1),
		(drawing, 1367, 1367, 0, 0, 0, 0, 1, 1),
		(drawing, 1366, 1366, 0, 0, 0, 0, 1, 1),
		(drawing, 1365, 1365, 0, 0, 0, 0, 1, 1),
		(drawing, 1364, 1364, 0, 0, 0, 0, 1, 1),
		(drawing, 1363, 1363, 0, 0, 0, 0, 1, 1),
		(drawing, 1362, 1362, 0, 0, 0, 0, 1, 1),
		(drawing, 1361, 1361, 0, 0, 0, 0, 1, 1),
		(drawing, 1360, 1360, 0, 0, 0, 0, 1, 1),
		(drawing, 1359, 1359, 0, 0, 0, 0, 1, 1),
		(drawing, 1358, 1358, 0, 0, 0, 0, 1, 1),
		(drawing, 1357, 1357, 0, 0, 0, 0, 1, 1),
		(drawing, 1356, 1356, 0, 0, 0, 0, 1, 1),
		(drawing, 1355, 1355, 0, 0, 0, 0, 1, 1),
		(drawing, 1354, 1354, 0, 0, 0, 0, 1, 1),
		(drawing, 1353, 1353, 0, 0, 0, 0, 1, 1),
		(drawing, 1352, 1352, 0, 0, 0, 0, 1, 1),
		(drawing, 1351, 1351, 0, 0, 0, 0, 1, 1),
		(drawing, 1350, 1350, 0, 0, 0, 0, 1, 1),
		(drawing, 1349, 1349, 0, 0, 0, 0, 1, 1),
		(drawing, 1348, 1348, 0, 0, 0, 0, 1, 1),
		(drawing, 1347, 1347, 0, 0, 0, 0, 1, 1),
		(drawing, 1346, 1346, 0, 0, 0, 0, 1, 1),
		(drawing, 1345, 1345, 0, 0, 0, 0, 1, 1),
		(drawing, 1344, 1344, 0, 0, 0, 0, 1, 1),
		(drawing, 1343, 1343, 0, 0, 0, 0, 1, 1),
		(drawing, 1342, 1342, 0, 0, 0, 0, 1, 1),
		(drawing, 1341, 1341, 0, 0, 0, 0, 1, 1),
		(drawing, 1340, 1340, 0, 0, 0, 0, 1, 1),
		(drawing, 1339, 1339, 0, 0, 0, 0, 1, 1),
		(drawing, 1338, 1338, 0, 0, 0, 0, 1, 1),
		(drawing, 1337, 1337, 0, 0, 0, 0, 1, 1),
		(drawing, 1336, 1336, 0, 0, 0, 0, 1, 1),
		(drawing, 1335, 1335, 0, 0, 0, 0, 1, 1),
		(drawing, 1334, 1334, 0, 0, 0, 0, 1, 1),
		(drawing, 1333, 1333, 0, 0, 0, 0, 1, 1),
		(drawing, 1332, 1332, 0, 0, 0, 0, 1, 1),
		(drawing, 1331, 1331, 0, 0, 0, 0, 1, 1),
		(drawing, 1330, 1330, 0, 0, 0, 0, 1, 1),
		(drawing, 1329, 1329, 0, 0, 0, 0, 1, 1),
		(drawing, 1328, 1328, 0, 0, 0, 0, 1, 1),
		(drawing, 1327, 1327, 0, 0, 0, 0, 1, 1),
		(drawing, 1326, 1326, 0, 0, 0, 0, 1, 1),
		(drawing, 1325, 1325, 0, 0, 0, 0, 1, 1),
		(drawing, 1324, 1324, 0, 0, 0, 0, 1, 1),
		(drawing, 1323, 1323, 0, 0, 0, 0, 1, 1),
		(drawing, 1322, 1322, 0, 0, 0, 0, 1, 1),
		(drawing, 1321, 1321, 0, 0, 0, 0, 1, 1),
		(drawing, 1320, 1320, 0, 0, 0, 0, 1, 1),
		(drawing, 1319, 1319, 0, 0, 0, 0, 1, 1),
		(drawing, 1318, 1318, 0, 0, 0, 0, 1, 1),
		(drawing, 1317, 1317, 0, 0, 0, 0, 1, 1),
		(drawing, 1316, 1316, 0, 0, 0, 0, 1, 1),
		(drawing, 1315, 1315, 0, 0, 0, 0, 1, 1),
		(drawing, 1314, 1314, 0, 0, 0, 0, 1, 1),
		(drawing, 1313, 1313, 0, 0, 0, 0, 1, 1),
		(drawing, 1312, 1312, 0, 0, 0, 0, 1, 1),
		(drawing, 1311, 1311, 0, 0, 0, 0, 1, 1),
		(drawing, 1310, 1310, 0, 0, 0, 0, 1, 1),
		(drawing, 1309, 1309, 0, 0, 0, 0, 1, 1),
		(drawing, 1308, 1308, 0, 0, 0, 0, 1, 1),
		(drawing, 1307, 1307, 0, 0, 0, 0, 1, 1),
		(drawing, 1306, 1306, 0, 0, 0, 0, 1, 1),
		(drawing, 1305, 1305, 0, 0, 0, 0, 1, 1),
		(drawing, 1304, 1304, 0, 0, 0, 0, 1, 1),
		(drawing, 1303, 1303, 0, 0, 0, 0, 1, 1),
		(drawing, 1302, 1302, 0, 0, 0, 0, 1, 1),
		(drawing, 1301, 1301, 0, 0, 0, 0, 1, 1),
		(drawing, 1300, 1300, 0, 0, 0, 0, 1, 1),
		(drawing, 1299, 1299, 0, 0, 0, 0, 1, 1),
		(drawing, 1298, 1298, 0, 0, 0, 0, 1, 1),
		(drawing, 1297, 1297, 0, 0, 0, 0, 1, 1),
		(drawing, 1296, 1296, 0, 0, 0, 0, 1, 1),
		(drawing, 1295, 1295, 0, 0, 0, 0, 1, 1),
		(drawing, 1294, 1294, 0, 0, 0, 0, 1, 1),
		(drawing, 1293, 1293, 0, 0, 0, 0, 1, 1),
		(drawing, 1292, 1292, 0, 0, 0, 0, 1, 1),
		(drawing, 1291, 1291, 0, 0, 0, 0, 1, 1),
		(drawing, 1290, 1290, 0, 0, 0, 0, 1, 1),
		(drawing, 1289, 1289, 0, 0, 0, 0, 1, 1),
		(drawing, 1288, 1288, 0, 0, 0, 0, 1, 1),
		(drawing, 1287, 1287, 0, 0, 0, 0, 1, 1),
		(drawing, 1286, 1286, 0, 0, 0, 0, 1, 1),
		(drawing, 1285, 1285, 0, 0, 0, 0, 1, 1),
		(drawing, 1284, 1284, 0, 0, 0, 0, 1, 1),
		(drawing, 1283, 1283, 0, 0, 0, 0, 1, 1),
		(drawing, 1282, 1282, 0, 0, 0, 0, 1, 1),
		(drawing, 1281, 1281, 0, 0, 0, 0, 1, 1),
		(drawing, 1280, 1280, 0, 0, 0, 0, 1, 1),
		(drawing, 1279, 1279, 0, 0, 0, 0, 1, 1),
		(drawing, 1278, 1278, 0, 0, 0, 0, 1, 1),
		(drawing, 1277, 1277, 0, 0, 0, 0, 1, 1),
		(drawing, 1276, 1276, 0, 0, 0, 0, 1, 1),
		(drawing, 1275, 1275, 0, 0, 0, 0, 1, 1),
		(drawing, 1274, 1274, 0, 0, 0, 0, 1, 1),
		(drawing, 1273, 1273, 0, 0, 0, 0, 1, 1),
		(drawing, 1272, 1272, 0, 0, 0, 0, 1, 1),
		(drawing, 1271, 1271, 0, 0, 0, 0, 1, 1),
		(drawing, 1270, 1270, 0, 0, 0, 0, 1, 1),
		(drawing, 1269, 1269, 0, 0, 0, 0, 1, 1),
		(drawing, 1268, 1268, 0, 0, 0, 0, 1, 1),
		(drawing, 1267, 1267, 0, 0, 0, 0, 1, 1),
		(drawing, 1266, 1266, 0, 0, 0, 0, 1, 1),
		(drawing, 1265, 1265, 0, 0, 0, 0, 1, 1),
		(drawing, 1264, 1264, 0, 0, 0, 0, 1, 1),
		(drawing, 1263, 1263, 0, 0, 0, 0, 1, 1),
		(drawing, 1262, 1262, 0, 0, 0, 0, 1, 1),
		(drawing, 1261, 1261, 0, 0, 0, 0, 1, 1),
		(drawing, 1260, 1260, 0, 0, 0, 0, 1, 1),
		(drawing, 1259, 1259, 0, 0, 0, 0, 1, 1),
		(drawing, 1258, 1258, 0, 0, 0, 0, 1, 1),
		(drawing, 1257, 1257, 0, 0, 0, 0, 1, 1),
		(drawing, 1256, 1256, 0, 0, 0, 0, 1, 1),
		(drawing, 1255, 1255, 0, 0, 0, 0, 1, 1),
		(drawing, 1254, 1254, 0, 0, 0, 0, 1, 1),
		(drawing, 1253, 1253, 0, 0, 0, 0, 1, 1),
		(drawing, 1252, 1252, 0, 0, 0, 0, 1, 1),
		(drawing, 1251, 1251, 0, 0, 0, 0, 1, 1),
		(drawing, 1250, 1250, 0, 0, 0, 0, 1, 1),
		(drawing, 1249, 1249, 0, 0, 0, 0, 1, 1),
		(drawing, 1248, 1248, 0, 0, 0, 0, 1, 1),
		(drawing, 1247, 1247, 0, 0, 0, 0, 1, 1),
		(drawing, 1246, 1246, 0, 0, 0, 0, 1, 1),
		(drawing, 1245, 1245, 0, 0, 0, 0, 1, 1),
		(drawing, 1244, 1244, 0, 0, 0, 0, 1, 1),
		(drawing, 1243, 1243, 0, 0, 0, 0, 1, 1),
		(drawing, 1242, 1242, 0, 0, 0, 0, 1, 1),
		(drawing, 1241, 1241, 0, 0, 0, 0, 1, 1),
		(drawing, 1240, 1240, 0, 0, 0, 0, 1, 1),
		(drawing, 1239, 1239, 0, 0, 0, 0, 1, 1),
		(drawing, 1238, 1238, 0, 0, 0, 0, 1, 1),
		(drawing, 1237, 1237, 0, 0, 0, 0, 1, 1),
		(drawing, 1236, 1236, 0, 0, 0, 0, 1, 1),
		(drawing, 1235, 1235, 0, 0, 0, 0, 1, 1),
		(drawing, 1234, 1234, 0, 0, 0, 0, 1, 1),
		(drawing, 1233, 1233, 0, 0, 0, 0, 1, 1),
		(drawing, 1232, 1232, 0, 0, 0, 0, 1, 1),
		(drawing, 1231, 1231, 0, 0, 0, 0, 1, 1),
		(drawing, 1230, 1230, 0, 0, 0, 0, 1, 1),
		(drawing, 1229, 1229, 0, 0, 0, 0, 1, 1),
		(drawing, 1228, 1228, 0, 0, 0, 0, 1, 1),
		(drawing, 1227, 1227, 0, 0, 0, 0, 1, 1),
		(drawing, 1226, 1226, 0, 0, 0, 0, 1, 1),
		(drawing, 1225, 1225, 0, 0, 0, 0, 1, 1),
		(drawing, 1224, 1224, 0, 0, 0, 0, 1, 1),
		(drawing, 1223, 1223, 0, 0, 0, 0, 1, 1),
		(drawing, 1222, 1222, 0, 0, 0, 0, 1, 1),
		(drawing, 1221, 1221, 0, 0, 0, 0, 1, 1),
		(drawing, 1220, 1220, 0, 0, 0, 0, 1, 1),
		(drawing, 1219, 1219, 0, 0, 0, 0, 1, 1),
		(drawing, 1218, 1218, 0, 0, 0, 0, 1, 1),
		(drawing, 1217, 1217, 0, 0, 0, 0, 1, 1),
		(drawing, 1216, 1216, 0, 0, 0, 0, 1, 1),
		(drawing, 1215, 1215, 0, 0, 0, 0, 1, 1),
		(drawing, 1214, 1214, 0, 0, 0, 0, 1, 1),
		(drawing, 1213, 1213, 0, 0, 0, 0, 1, 1),
		(drawing, 1212, 1212, 0, 0, 0, 0, 1, 1),
		(drawing, 1211, 1211, 0, 0, 0, 0, 1, 1),
		(drawing, 1210, 1210, 0, 0, 0, 0, 1, 1),
		(drawing, 1209, 1209, 0, 0, 0, 0, 1, 1),
		(drawing, 1208, 1208, 0, 0, 0, 0, 1, 1),
		(drawing, 1207, 1207, 0, 0, 0, 0, 1, 1),
		(drawing, 1206, 1206, 0, 0, 0, 0, 1, 1),
		(drawing, 1205, 1205, 0, 0, 0, 0, 1, 1),
		(drawing, 1204, 1204, 0, 0, 0, 0, 1, 1),
		(drawing, 1203, 1203, 0, 0, 0, 0, 1, 1),
		(drawing, 1202, 1202, 0, 0, 0, 0, 1, 1),
		(drawing, 1201, 1201, 0, 0, 0, 0, 1, 1),
		(drawing, 1200, 1200, 0, 0, 0, 0, 1, 1),
		(drawing, 1199, 1199, 0, 0, 0, 0, 1, 1),
		(drawing, 1198, 1198, 0, 0, 0, 0, 1, 1),
		(drawing, 1197, 1197, 0, 0, 0, 0, 1, 1),
		(drawing, 1196, 1196, 0, 0, 0, 0, 1, 1),
		(drawing, 1195, 1195, 0, 0, 0, 0, 1, 1),
		(drawing, 1194, 1194, 0, 0, 0, 0, 1, 1),
		(drawing, 1193, 1193, 0, 0, 0, 0, 1, 1),
		(drawing, 1192, 1192, 0, 0, 0, 0, 1, 1),
		(drawing, 1191, 1191, 0, 0, 0, 0, 1, 1),
		(drawing, 1190, 1190, 0, 0, 0, 0, 1, 1),
		(drawing, 1189, 1189, 0, 0, 0, 0, 1, 1),
		(drawing, 1188, 1188, 0, 0, 0, 0, 1, 1),
		(drawing, 1187, 1187, 0, 0, 0, 0, 1, 1),
		(drawing, 1186, 1186, 0, 0, 0, 0, 1, 1),
		(drawing, 1185, 1185, 0, 0, 0, 0, 1, 1),
		(drawing, 1184, 1184, 0, 0, 0, 0, 1, 1),
		(drawing, 1183, 1183, 0, 0, 0, 0, 1, 1),
		(drawing, 1182, 1182, 0, 0, 0, 0, 1, 1),
		(drawing, 1181, 1181, 0, 0, 0, 0, 1, 1),
		(drawing, 1180, 1180, 0, 0, 0, 0, 1, 1),
		(drawing, 1179, 1179, 0, 0, 0, 0, 1, 1),
		(drawing, 1178, 1178, 0, 0, 0, 0, 1, 1),
		(drawing, 1177, 1177, 0, 0, 0, 0, 1, 1),
		(drawing, 1176, 1176, 0, 0, 0, 0, 1, 1),
		(drawing, 1175, 1175, 0, 0, 0, 0, 1, 1),
		(drawing, 1174, 1174, 0, 0, 0, 0, 1, 1),
		(drawing, 1173, 1173, 0, 0, 0, 0, 1, 1),
		(drawing, 1172, 1172, 0, 0, 0, 0, 1, 1),
		(drawing, 1171, 1171, 0, 0, 0, 0, 1, 1),
		(drawing, 1170, 1170, 0, 0, 0, 0, 1, 1),
		(drawing, 1169, 1169, 0, 0, 0, 0, 1, 1),
		(drawing, 1168, 1168, 0, 0, 0, 0, 1, 1),
		(drawing, 1167, 1167, 0, 0, 0, 0, 1, 1),
		(drawing, 1166, 1166, 0, 0, 0, 0, 1, 1),
		(drawing, 1165, 1165, 0, 0, 0, 0, 1, 1),
		(drawing, 1164, 1164, 0, 0, 0, 0, 1, 1),
		(drawing, 1163, 1163, 0, 0, 0, 0, 1, 1),
		(drawing, 1162, 1162, 0, 0, 0, 0, 1, 1),
		(drawing, 1161, 1161, 0, 0, 0, 0, 1, 1),
		(drawing, 1160, 1160, 0, 0, 0, 0, 1, 1),
		(drawing, 1159, 1159, 0, 0, 0, 0, 1, 1),
		(drawing, 1158, 1158, 0, 0, 0, 0, 1, 1),
		(drawing, 1157, 1157, 0, 0, 0, 0, 1, 1),
		(drawing, 1156, 1156, 0, 0, 0, 0, 1, 1),
		(drawing, 1155, 1155, 0, 0, 0, 0, 1, 1),
		(drawing, 1154, 1154, 0, 0, 0, 0, 1, 1),
		(drawing, 1153, 1153, 0, 0, 0, 0, 1, 1),
		(drawing, 1152, 1152, 0, 0, 0, 0, 1, 1),
		(drawing, 1151, 1151, 0, 0, 0, 0, 1, 1),
		(drawing, 1150, 1150, 0, 0, 0, 0, 1, 1),
		(drawing, 1149, 1149, 0, 0, 0, 0, 1, 1),
		(drawing, 1148, 1148, 0, 0, 0, 0, 1, 1),
		(drawing, 1147, 1147, 0, 0, 0, 0, 1, 1),
		(drawing, 1146, 1146, 0, 0, 0, 0, 1, 1),
		(drawing, 1145, 1145, 0, 0, 0, 0, 1, 1),
		(drawing, 1144, 1144, 0, 0, 0, 0, 1, 1),
		(drawing, 1143, 1143, 0, 0, 0, 0, 1, 1),
		(drawing, 1142, 1142, 0, 0, 0, 0, 1, 1),
		(drawing, 1141, 1141, 0, 0, 0, 0, 1, 1),
		(drawing, 1140, 1140, 0, 0, 0, 0, 1, 1),
		(drawing, 1139, 1139, 0, 0, 0, 0, 1, 1),
		(drawing, 1138, 1138, 0, 0, 0, 0, 1, 1),
		(drawing, 1137, 1137, 0, 0, 0, 0, 1, 1),
		(drawing, 1136, 1136, 0, 0, 0, 0, 1, 1),
		(drawing, 1135, 1135, 0, 0, 0, 0, 1, 1),
		(drawing, 1134, 1134, 0, 0, 0, 0, 1, 1),
		(drawing, 1133, 1133, 0, 0, 0, 0, 1, 1),
		(drawing, 1132, 1132, 0, 0, 0, 0, 1, 1),
		(drawing, 1131, 1131, 0, 0, 0, 0, 1, 1),
		(drawing, 1130, 1130, 0, 0, 0, 0, 1, 1),
		(drawing, 1129, 1129, 0, 0, 0, 0, 1, 1),
		(drawing, 1128, 1128, 0, 0, 0, 0, 1, 1),
		(drawing, 1127, 1127, 0, 0, 0, 0, 1, 1),
		(drawing, 1126, 1126, 0, 0, 0, 0, 1, 1),
		(drawing, 1125, 1125, 0, 0, 0, 0, 1, 1),
		(drawing, 1124, 1124, 0, 0, 0, 0, 1, 1),
		(drawing, 1123, 1123, 0, 0, 0, 0, 1, 1),
		(drawing, 1122, 1122, 0, 0, 0, 0, 1, 1),
		(drawing, 1121, 1121, 0, 0, 0, 0, 1, 1),
		(drawing, 1120, 1120, 0, 0, 0, 0, 1, 1),
		(drawing, 1119, 1119, 0, 0, 0, 0, 1, 1),
		(drawing, 1118, 1118, 0, 0, 0, 0, 1, 1),
		(drawing, 1117, 1117, 0, 0, 0, 0, 1, 1),
		(drawing, 1116, 1116, 0, 0, 0, 0, 1, 1),
		(drawing, 1115, 1115, 0, 0, 0, 0, 1, 1),
		(drawing, 1114, 1114, 0, 0, 0, 0, 1, 1),
		(drawing, 1113, 1113, 0, 0, 0, 0, 1, 1),
		(drawing, 1112, 1112, 0, 0, 0, 0, 1, 1),
		(drawing, 1111, 1111, 0, 0, 0, 0, 1, 1),
		(drawing, 1110, 1110, 0, 0, 0, 0, 1, 1),
		(drawing, 1109, 1109, 0, 0, 0, 0, 1, 1),
		(drawing, 1108, 1108, 0, 0, 0, 0, 1, 1),
		(drawing, 1107, 1107, 0, 0, 0, 0, 1, 1),
		(drawing, 1106, 1106, 0, 0, 0, 0, 1, 1),
		(drawing, 1105, 1105, 0, 0, 0, 0, 1, 1),
		(drawing, 1104, 1104, 0, 0, 0, 0, 1, 1),
		(drawing, 1103, 1103, 0, 0, 0, 0, 1, 1),
		(drawing, 1102, 1102, 0, 0, 0, 0, 1, 1),
		(drawing, 1101, 1101, 0, 0, 0, 0, 1, 1),
		(drawing, 1100, 1100, 0, 0, 0, 0, 1, 1),
		(drawing, 1099, 1099, 0, 0, 0, 0, 1, 1),
		(drawing, 1098, 1098, 0, 0, 0, 0, 1, 1),
		(drawing, 1097, 1097, 0, 0, 0, 0, 1, 1),
		(drawing, 1096, 1096, 0, 0, 0, 0, 1, 1),
		(drawing, 1095, 1095, 0, 0, 0, 0, 1, 1),
		(drawing, 1094, 1094, 0, 0, 0, 0, 1, 1),
		(drawing, 1093, 1093, 0, 0, 0, 0, 1, 1),
		(drawing, 1092, 1092, 0, 0, 0, 0, 1, 1),
		(drawing, 1091, 1091, 0, 0, 0, 0, 1, 1),
		(drawing, 1090, 1090, 0, 0, 0, 0, 1, 1),
		(drawing, 1089, 1089, 0, 0, 0, 0, 1, 1),
		(drawing, 1088, 1088, 0, 0, 0, 0, 1, 1),
		(drawing, 1087, 1087, 0, 0, 0, 0, 1, 1),
		(drawing, 1086, 1086, 0, 0, 0, 0, 1, 1),
		(drawing, 1085, 1085, 0, 0, 0, 0, 1, 1),
		(drawing, 1084, 1084, 0, 0, 0, 0, 1, 1),
		(drawing, 1083, 1083, 0, 0, 0, 0, 1, 1),
		(drawing, 1082, 1082, 0, 0, 0, 0, 1, 1),
		(drawing, 1081, 1081, 0, 0, 0, 0, 1, 1),
		(drawing, 1080, 1080, 0, 0, 0, 0, 1, 1),
		(drawing, 1079, 1079, 0, 0, 0, 0, 1, 1),
		(drawing, 1078, 1078, 0, 0, 0, 0, 1, 1),
		(drawing, 1077, 1077, 0, 0, 0, 0, 1, 1),
		(drawing, 1076, 1076, 0, 0, 0, 0, 1, 1),
		(drawing, 1075, 1075, 0, 0, 0, 0, 1, 1),
		(drawing, 1074, 1074, 0, 0, 0, 0, 1, 1),
		(drawing, 1073, 1073, 0, 0, 0, 0, 1, 1),
		(drawing, 1072, 1072, 0, 0, 0, 0, 1, 1),
		(drawing, 1071, 1071, 0, 0, 0, 0, 1, 1),
		(drawing, 1070, 1070, 0, 0, 0, 0, 1, 1),
		(drawing, 1069, 1069, 0, 0, 0, 0, 1, 1),
		(drawing, 1068, 1068, 0, 0, 0, 0, 1, 1),
		(drawing, 1067, 1067, 0, 0, 0, 0, 1, 1),
		(drawing, 1066, 1066, 0, 0, 0, 0, 1, 1),
		(drawing, 1065, 1065, 0, 0, 0, 0, 1, 1),
		(drawing, 1064, 1064, 0, 0, 0, 0, 1, 1),
		(drawing, 1063, 1063, 0, 0, 0, 0, 1, 1),
		(drawing, 1062, 1062, 0, 0, 0, 0, 1, 1),
		(drawing, 1061, 1061, 0, 0, 0, 0, 1, 1),
		(drawing, 1060, 1060, 0, 0, 0, 0, 1, 1),
		(drawing, 1059, 1059, 0, 0, 0, 0, 1, 1),
		(drawing, 1058, 1058, 0, 0, 0, 0, 1, 1),
		(drawing, 1057, 1057, 0, 0, 0, 0, 1, 1),
		(drawing, 1056, 1056, 0, 0, 0, 0, 1, 1),
		(drawing, 1055, 1055, 0, 0, 0, 0, 1, 1),
		(drawing, 1054, 1054, 0, 0, 0, 0, 1, 1),
		(drawing, 1053, 1053, 0, 0, 0, 0, 1, 1),
		(drawing, 1052, 1052, 0, 0, 0, 0, 1, 1),
		(drawing, 1051, 1051, 0, 0, 0, 0, 1, 1),
		(drawing, 1050, 1050, 0, 0, 0, 0, 1, 1),
		(drawing, 1049, 1049, 0, 0, 0, 0, 1, 1),
		(drawing, 1048, 1048, 0, 0, 0, 0, 1, 1),
		(drawing, 1047, 1047, 0, 0, 0, 0, 1, 1),
		(drawing, 1046, 1046, 0, 0, 0, 0, 1, 1),
		(drawing, 1045, 1045, 0, 0, 0, 0, 1, 1),
		(drawing, 1044, 1044, 0, 0, 0, 0, 1, 1),
		(drawing, 1043, 1043, 0, 0, 0, 0, 1, 1),
		(drawing, 1042, 1042, 0, 0, 0, 0, 1, 1),
		(drawing, 1041, 1041, 0, 0, 0, 0, 1, 1),
		(drawing, 1040, 1040, 0, 0, 0, 0, 1, 1),
		(drawing, 1039, 1039, 0, 0, 0, 0, 1, 1),
		(drawing, 1038, 1038, 0, 0, 0, 0, 1, 1),
		(drawing, 1037, 1037, 0, 0, 0, 0, 1, 1),
		(drawing, 1036, 1036, 0, 0, 0, 0, 1, 1),
		(drawing, 1035, 1035, 0, 0, 0, 0, 1, 1),
		(drawing, 1034, 1034, 0, 0, 0, 0, 1, 1),
		(drawing, 1033, 1033, 0, 0, 0, 0, 1, 1),
		(drawing, 1032, 1032, 0, 0, 0, 0, 1, 1),
		(drawing, 1031, 1031, 0, 0, 0, 0, 1, 1),
		(drawing, 1030, 1030, 0, 0, 0, 0, 1, 1),
		(drawing, 1029, 1029, 0, 0, 0, 0, 1, 1),
		(drawing, 1028, 1028, 0, 0, 0, 0, 1, 1),
		(drawing, 1027, 1027, 0, 0, 0, 0, 1, 1),
		(drawing, 1026, 1026, 0, 0, 0, 0, 1, 1),
		(drawing, 1025, 1025, 0, 0, 0, 0, 1, 1),
		(drawing, 1024, 1024, 0, 0, 0, 0, 1, 1),
		(drawing, 1023, 1023, 0, 0, 0, 0, 1, 1),
		(drawing, 1022, 1022, 0, 0, 0, 0, 1, 1),
		(drawing, 1021, 1021, 0, 0, 0, 0, 1, 1),
		(drawing, 1020, 1020, 0, 0, 0, 0, 1, 1),
		(drawing, 1019, 1019, 0, 0, 0, 0, 1, 1),
		(drawing, 1018, 1018, 0, 0, 0, 0, 1, 1),
		(drawing, 1017, 1017, 0, 0, 0, 0, 1, 1),
		(drawing, 1016, 1016, 0, 0, 0, 0, 1, 1),
		(drawing, 1015, 1015, 0, 0, 0, 0, 1, 1),
		(drawing, 1014, 1014, 0, 0, 0, 0, 1, 1),
		(drawing, 1013, 1013, 0, 0, 0, 0, 1, 1),
		(drawing, 1012, 1012, 0, 0, 0, 0, 1, 1),
		(drawing, 1011, 1011, 0, 0, 0, 0, 1, 1),
		(drawing, 1010, 1010, 0, 0, 0, 0, 1, 1),
		(drawing, 1009, 1009, 0, 0, 0, 0, 1, 1),
		(drawing, 1008, 1008, 0, 0, 0, 0, 1, 1),
		(drawing, 1007, 1007, 0, 0, 0, 0, 1, 1),
		(drawing, 1006, 1006, 0, 0, 0, 0, 1, 1),
		(drawing, 1005, 1005, 0, 0, 0, 0, 1, 1),
		(drawing, 1004, 1004, 0, 0, 0, 0, 1, 1),
		(drawing, 1003, 1003, 0, 0, 0, 0, 1, 1),
		(drawing, 1002, 1002, 0, 0, 0, 0, 1, 1),
		(drawing, 1001, 1001, 0, 0, 0, 0, 1, 1),
		(drawing, 1000, 1000, 0, 0, 0, 0, 1, 1),
		(drawing, 999, 999, 0, 0, 0, 0, 1, 1),
		(drawing, 998, 998, 0, 0, 0, 0, 1, 1),
		(drawing, 997, 997, 0, 0, 0, 0, 1, 1),
		(drawing, 996, 996, 0, 0, 0, 0, 1, 1),
		(drawing, 995, 995, 0, 0, 0, 0, 1, 1),
		(drawing, 994, 994, 0, 0, 0, 0, 1, 1),
		(drawing, 993, 993, 0, 0, 0, 0, 1, 1),
		(drawing, 992, 992, 0, 0, 0, 0, 1, 1),
		(drawing, 991, 991, 0, 0, 0, 0, 1, 1),
		(drawing, 990, 990, 0, 0, 0, 0, 1, 1),
		(drawing, 989, 989, 0, 0, 0, 0, 1, 1),
		(drawing, 988, 988, 0, 0, 0, 0, 1, 1),
		(drawing, 987, 987, 0, 0, 0, 0, 1, 1),
		(drawing, 986, 986, 0, 0, 0, 0, 1, 1),
		(drawing, 985, 985, 0, 0, 0, 0, 1, 1),
		(drawing, 984, 984, 0, 0, 0, 0, 1, 1),
		(drawing, 983, 983, 0, 0, 0, 0, 1, 1),
		(drawing, 982, 982, 0, 0, 0, 0, 1, 1),
		(drawing, 981, 981, 0, 0, 0, 0, 1, 1),
		(drawing, 980, 980, 0, 0, 0, 0, 1, 1),
		(drawing, 979, 979, 0, 0, 0, 0, 1, 1),
		(drawing, 978, 978, 0, 0, 0, 0, 1, 1),
		(drawing, 977, 977, 0, 0, 0, 0, 1, 1),
		(drawing, 976, 976, 0, 0, 0, 0, 1, 1),
		(drawing, 975, 975, 0, 0, 0, 0, 1, 1),
		(drawing, 974, 974, 0, 0, 0, 0, 1, 1),
		(drawing, 973, 973, 0, 0, 0, 0, 1, 1),
		(drawing, 972, 972, 0, 0, 0, 0, 1, 1),
		(drawing, 971, 971, 0, 0, 0, 0, 1, 1),
		(drawing, 970, 970, 0, 0, 0, 0, 1, 1),
		(drawing, 969, 969, 0, 0, 0, 0, 1, 1),
		(drawing, 968, 968, 0, 0, 0, 0, 1, 1),
		(drawing, 967, 967, 0, 0, 0, 0, 1, 1),
		(drawing, 966, 966, 0, 0, 0, 0, 1, 1),
		(drawing, 965, 965, 0, 0, 0, 0, 1, 1),
		(drawing, 964, 964, 0, 0, 0, 0, 1, 1),
		(drawing, 963, 963, 0, 0, 0, 0, 1, 1),
		(drawing, 962, 962, 0, 0, 0, 0, 1, 1),
		(drawing, 961, 961, 0, 0, 0, 0, 1, 1),
		(drawing, 960, 960, 0, 0, 0, 0, 1, 1),
		(drawing, 959, 959, 0, 0, 0, 0, 1, 1),
		(drawing, 958, 958, 0, 0, 0, 0, 1, 1),
		(drawing, 957, 957, 0, 0, 0, 0, 1, 1),
		(drawing, 956, 956, 0, 0, 0, 0, 1, 1),
		(drawing, 955, 955, 0, 0, 0, 0, 1, 1),
		(drawing, 954, 954, 0, 0, 0, 0, 1, 1),
		(drawing, 953, 953, 0, 0, 0, 0, 1, 1),
		(drawing, 952, 952, 0, 0, 0, 0, 1, 1),
		(drawing, 951, 951, 0, 0, 0, 0, 1, 1),
		(drawing, 950, 950, 0, 0, 0, 0, 1, 1),
		(drawing, 949, 949, 0, 0, 0, 0, 1, 1),
		(drawing, 948, 948, 0, 0, 0, 0, 1, 1),
		(drawing, 947, 947, 0, 0, 0, 0, 1, 1),
		(drawing, 946, 946, 0, 0, 0, 0, 1, 1),
		(drawing, 945, 945, 0, 0, 0, 0, 1, 1),
		(drawing, 944, 944, 0, 0, 0, 0, 1, 1),
		(drawing, 943, 943, 0, 0, 0, 0, 1, 1),
		(drawing, 942, 942, 0, 0, 0, 0, 1, 1),
		(drawing, 941, 941, 0, 0, 0, 0, 1, 1),
		(drawing, 940, 940, 0, 0, 0, 0, 1, 1),
		(drawing, 939, 939, 0, 0, 0, 0, 1, 1),
		(drawing, 938, 938, 0, 0, 0, 0, 1, 1),
		(drawing, 937, 937, 0, 0, 0, 0, 1, 1),
		(drawing, 936, 936, 0, 0, 0, 0, 1, 1),
		(drawing, 935, 935, 0, 0, 0, 0, 1, 1),
		(drawing, 934, 934, 0, 0, 0, 0, 1, 1),
		(drawing, 933, 933, 0, 0, 0, 0, 1, 1),
		(drawing, 932, 932, 0, 0, 0, 0, 1, 1),
		(drawing, 931, 931, 0, 0, 0, 0, 1, 1),
		(drawing, 930, 930, 0, 0, 0, 0, 1, 1),
		(drawing, 929, 929, 0, 0, 0, 0, 1, 1),
		(drawing, 928, 928, 0, 0, 0, 0, 1, 1),
		(drawing, 927, 927, 0, 0, 0, 0, 1, 1),
		(drawing, 926, 926, 0, 0, 0, 0, 1, 1),
		(drawing, 925, 925, 0, 0, 0, 0, 1, 1),
		(drawing, 924, 924, 0, 0, 0, 0, 1, 1),
		(drawing, 923, 923, 0, 0, 0, 0, 1, 1),
		(drawing, 922, 922, 0, 0, 0, 0, 1, 1),
		(drawing, 921, 921, 0, 0, 0, 0, 1, 1),
		(drawing, 920, 920, 0, 0, 0, 0, 1, 1),
		(drawing, 919, 919, 0, 0, 0, 0, 1, 1),
		(drawing, 918, 918, 0, 0, 0, 0, 1, 1),
		(drawing, 917, 917, 0, 0, 0, 0, 1, 1),
		(drawing, 916, 916, 0, 0, 0, 0, 1, 1),
		(drawing, 915, 915, 0, 0, 0, 0, 1, 1),
		(drawing, 914, 914, 0, 0, 0, 0, 1, 1),
		(drawing, 913, 913, 0, 0, 0, 0, 1, 1),
		(drawing, 912, 912, 0, 0, 0, 0, 1, 1),
		(drawing, 911, 911, 0, 0, 0, 0, 1, 1),
		(drawing, 910, 910, 0, 0, 0, 0, 1, 1),
		(drawing, 909, 909, 0, 0, 0, 0, 1, 1),
		(drawing, 908, 908, 0, 0, 0, 0, 1, 1),
		(drawing, 907, 907, 0, 0, 0, 0, 1, 1),
		(drawing, 906, 906, 0, 0, 0, 0, 1, 1),
		(drawing, 905, 905, 0, 0, 0, 0, 1, 1),
		(drawing, 904, 904, 0, 0, 0, 0, 1, 1),
		(drawing, 903, 903, 0, 0, 0, 0, 1, 1),
		(drawing, 902, 902, 0, 0, 0, 0, 1, 1),
		(drawing, 901, 901, 0, 0, 0, 0, 1, 1),
		(drawing, 900, 900, 0, 0, 0, 0, 1, 1),
		(drawing, 899, 899, 0, 0, 0, 0, 1, 1),
		(drawing, 898, 898, 0, 0, 0, 0, 1, 1),
		(drawing, 897, 897, 0, 0, 0, 0, 1, 1),
		(drawing, 896, 896, 0, 0, 0, 0, 1, 1),
		(drawing, 895, 895, 0, 0, 0, 0, 1, 1),
		(drawing, 894, 894, 0, 0, 0, 0, 1, 1),
		(drawing, 893, 893, 0, 0, 0, 0, 1, 1),
		(drawing, 892, 892, 0, 0, 0, 0, 1, 1),
		(drawing, 891, 891, 0, 0, 0, 0, 1, 1),
		(drawing, 890, 890, 0, 0, 0, 0, 1, 1),
		(drawing, 889, 889, 0, 0, 0, 0, 1, 1),
		(drawing, 888, 888, 0, 0, 0, 0, 1, 1),
		(drawing, 887, 887, 0, 0, 0, 0, 1, 1),
		(drawing, 886, 886, 0, 0, 0, 0, 1, 1),
		(drawing, 885, 885, 0, 0, 0, 0, 1, 1),
		(drawing, 884, 884, 0, 0, 0, 0, 1, 1),
		(drawing, 883, 883, 0, 0, 0, 0, 1, 1),
		(drawing, 882, 882, 0, 0, 0, 0, 1, 1),
		(drawing, 881, 881, 0, 0, 0, 0, 1, 1),
		(drawing, 880, 880, 0, 0, 0, 0, 1, 1),
		(drawing, 879, 879, 0, 0, 0, 0, 1, 1),
		(drawing, 878, 878, 0, 0, 0, 0, 1, 1),
		(drawing, 877, 877, 0, 0, 0, 0, 1, 1),
		(drawing, 876, 876, 0, 0, 0, 0, 1, 1),
		(drawing, 875, 875, 0, 0, 0, 0, 1, 1),
		(drawing, 874, 874, 0, 0, 0, 0, 1, 1),
		(drawing, 873, 873, 0, 0, 0, 0, 1, 1),
		(drawing, 872, 872, 0, 0, 0, 0, 1, 1),
		(drawing, 871, 871, 0, 0, 0, 0, 1, 1),
		(drawing, 870, 870, 0, 0, 0, 0, 1, 1),
		(drawing, 869, 869, 0, 0, 0, 0, 1, 1),
		(drawing, 868, 868, 0, 0, 0, 0, 1, 1),
		(drawing, 867, 867, 0, 0, 0, 0, 1, 1),
		(drawing, 866, 866, 0, 0, 0, 0, 1, 1),
		(drawing, 865, 865, 0, 0, 0, 0, 1, 1),
		(drawing, 864, 864, 0, 0, 0, 0, 1, 1),
		(drawing, 863, 863, 0, 0, 0, 0, 1, 1),
		(drawing, 862, 862, 0, 0, 0, 0, 1, 1),
		(drawing, 861, 861, 0, 0, 0, 0, 1, 1),
		(drawing, 860, 860, 0, 0, 0, 0, 1, 1),
		(drawing, 859, 859, 0, 0, 0, 0, 1, 1),
		(drawing, 858, 858, 0, 0, 0, 0, 1, 1),
		(drawing, 857, 857, 0, 0, 0, 0, 1, 1),
		(drawing, 856, 856, 0, 0, 0, 0, 1, 1),
		(drawing, 855, 855, 0, 0, 0, 0, 1, 1),
		(drawing, 854, 854, 0, 0, 0, 0, 1, 1),
		(drawing, 853, 853, 0, 0, 0, 0, 1, 1),
		(drawing, 852, 852, 0, 0, 0, 0, 1, 1),
		(drawing, 851, 851, 0, 0, 0, 0, 1, 1),
		(drawing, 850, 850, 0, 0, 0, 0, 1, 1),
		(drawing, 849, 849, 0, 0, 0, 0, 1, 1),
		(drawing, 848, 848, 0, 0, 0, 0, 1, 1),
		(drawing, 847, 847, 0, 0, 0, 0, 1, 1),
		(drawing, 846, 846, 0, 0, 0, 0, 1, 1),
		(drawing, 845, 845, 0, 0, 0, 0, 1, 1),
		(drawing, 844, 844, 0, 0, 0, 0, 1, 1),
		(drawing, 843, 843, 0, 0, 0, 0, 1, 1),
		(drawing, 842, 842, 0, 0, 0, 0, 1, 1),
		(drawing, 841, 841, 0, 0, 0, 0, 1, 1),
		(drawing, 840, 840, 0, 0, 0, 0, 1, 1),
		(drawing, 839, 839, 0, 0, 0, 0, 1, 1),
		(drawing, 838, 838, 0, 0, 0, 0, 1, 1),
		(drawing, 837, 837, 0, 0, 0, 0, 1, 1),
		(drawing, 836, 836, 0, 0, 0, 0, 1, 1),
		(drawing, 835, 835, 0, 0, 0, 0, 1, 1),
		(drawing, 834, 834, 0, 0, 0, 0, 1, 1),
		(drawing, 833, 833, 0, 0, 0, 0, 1, 1),
		(drawing, 832, 832, 0, 0, 0, 0, 1, 1),
		(drawing, 831, 831, 0, 0, 0, 0, 1, 1),
		(drawing, 830, 830, 0, 0, 0, 0, 1, 1),
		(drawing, 829, 829, 0, 0, 0, 0, 1, 1),
		(drawing, 828, 828, 0, 0, 0, 0, 1, 1),
		(drawing, 827, 827, 0, 0, 0, 0, 1, 1),
		(drawing, 826, 826, 0, 0, 0, 0, 1, 1),
		(drawing, 825, 825, 0, 0, 0, 0, 1, 1),
		(drawing, 824, 824, 0, 0, 0, 0, 1, 1),
		(drawing, 823, 823, 0, 0, 0, 0, 1, 1),
		(drawing, 822, 822, 0, 0, 0, 0, 1, 1),
		(drawing, 821, 821, 0, 0, 0, 0, 1, 1),
		(drawing, 820, 820, 0, 0, 0, 0, 1, 1),
		(drawing, 819, 819, 0, 0, 0, 0, 1, 1),
		(drawing, 818, 818, 0, 0, 0, 0, 1, 1),
		(drawing, 817, 817, 0, 0, 0, 0, 1, 1),
		(drawing, 816, 816, 0, 0, 0, 0, 1, 1),
		(drawing, 815, 815, 0, 0, 0, 0, 1, 1),
		(drawing, 814, 814, 0, 0, 0, 0, 1, 1),
		(drawing, 813, 813, 0, 0, 0, 0, 1, 1),
		(drawing, 812, 812, 0, 0, 0, 0, 1, 1),
		(drawing, 811, 811, 0, 0, 0, 0, 1, 1),
		(drawing, 810, 810, 0, 0, 0, 0, 1, 1),
		(drawing, 809, 809, 0, 0, 0, 0, 1, 1),
		(drawing, 808, 808, 0, 0, 0, 0, 1, 1),
		(drawing, 807, 807, 0, 0, 0, 0, 1, 1),
		(drawing, 806, 806, 0, 0, 0, 0, 1, 1),
		(drawing, 805, 805, 0, 0, 0, 0, 1, 1),
		(drawing, 804, 804, 0, 0, 0, 0, 1, 1),
		(drawing, 803, 803, 0, 0, 0, 0, 1, 1),
		(drawing, 802, 802, 0, 0, 0, 0, 1, 1),
		(drawing, 801, 801, 0, 0, 0, 0, 1, 1),
		(drawing, 800, 800, 0, 0, 0, 0, 1, 1),
		(drawing, 799, 799, 0, 0, 0, 0, 1, 1),
		(drawing, 798, 798, 0, 0, 0, 0, 1, 1),
		(drawing, 797, 797, 0, 0, 0, 0, 1, 1),
		(drawing, 796, 796, 0, 0, 0, 0, 1, 1),
		(drawing, 795, 795, 0, 0, 0, 0, 1, 1),
		(drawing, 794, 794, 0, 0, 0, 0, 1, 1),
		(drawing, 793, 793, 0, 0, 0, 0, 1, 1),
		(drawing, 792, 792, 0, 0, 0, 0, 1, 1),
		(drawing, 791, 791, 0, 0, 0, 0, 1, 1),
		(drawing, 790, 790, 0, 0, 0, 0, 1, 1),
		(drawing, 789, 789, 0, 0, 0, 0, 1, 1),
		(drawing, 788, 788, 0, 0, 0, 0, 1, 1),
		(drawing, 787, 787, 0, 0, 0, 0, 1, 1),
		(drawing, 786, 786, 0, 0, 0, 0, 1, 1),
		(drawing, 785, 785, 0, 0, 0, 0, 1, 1),
		(drawing, 784, 784, 0, 0, 0, 0, 1, 1),
		(drawing, 783, 783, 0, 0, 0, 0, 1, 1),
		(drawing, 782, 782, 0, 0, 0, 0, 1, 1),
		(drawing, 781, 781, 0, 0, 0, 0, 1, 1),
		(drawing, 780, 780, 0, 0, 0, 0, 1, 1),
		(drawing, 779, 779, 0, 0, 0, 0, 1, 1),
		(drawing, 778, 778, 0, 0, 0, 0, 1, 1),
		(drawing, 777, 777, 0, 0, 0, 0, 1, 1),
		(drawing, 776, 776, 0, 0, 0, 0, 1, 1),
		(drawing, 775, 775, 0, 0, 0, 0, 1, 1),
		(drawing, 774, 774, 0, 0, 0, 0, 1, 1),
		(drawing, 773, 773, 0, 0, 0, 0, 1, 1),
		(drawing, 772, 772, 0, 0, 0, 0, 1, 1),
		(drawing, 771, 771, 0, 0, 0, 0, 1, 1),
		(drawing, 770, 770, 0, 0, 0, 0, 1, 1),
		(drawing, 769, 769, 0, 0, 0, 0, 1, 1),
		(drawing, 768, 768, 0, 0, 0, 0, 1, 1),
		(drawing, 767, 767, 0, 0, 0, 0, 1, 1),
		(drawing, 766, 766, 0, 0, 0, 0, 1, 1),
		(drawing, 765, 765, 0, 0, 0, 0, 1, 1),
		(drawing, 764, 764, 0, 0, 0, 0, 1, 1),
		(drawing, 763, 763, 0, 0, 0, 0, 1, 1),
		(drawing, 762, 762, 0, 0, 0, 0, 1, 1),
		(drawing, 761, 761, 0, 0, 0, 0, 1, 1),
		(drawing, 760, 760, 0, 0, 0, 0, 1, 1),
		(drawing, 759, 759, 0, 0, 0, 0, 1, 1),
		(drawing, 758, 758, 0, 0, 0, 0, 1, 1),
		(drawing, 757, 757, 0, 0, 0, 0, 1, 1),
		(drawing, 756, 756, 0, 0, 0, 0, 1, 1),
		(drawing, 755, 755, 0, 0, 0, 0, 1, 1),
		(drawing, 754, 754, 0, 0, 0, 0, 1, 1),
		(drawing, 753, 753, 0, 0, 0, 0, 1, 1),
		(drawing, 752, 752, 0, 0, 0, 0, 1, 1),
		(drawing, 751, 751, 0, 0, 0, 0, 1, 1),
		(drawing, 750, 750, 0, 0, 0, 0, 1, 1),
		(drawing, 749, 749, 0, 0, 0, 0, 1, 1),
		(drawing, 748, 748, 0, 0, 0, 0, 1, 1),
		(drawing, 747, 747, 0, 0, 0, 0, 1, 1),
		(drawing, 746, 746, 0, 0, 0, 0, 1, 1),
		(drawing, 745, 745, 0, 0, 0, 0, 1, 1),
		(drawing, 744, 744, 0, 0, 0, 0, 1, 1),
		(drawing, 743, 743, 0, 0, 0, 0, 1, 1),
		(drawing, 742, 742, 0, 0, 0, 0, 1, 1),
		(drawing, 741, 741, 0, 0, 0, 0, 1, 1),
		(drawing, 740, 740, 0, 0, 0, 0, 1, 1),
		(drawing, 739, 739, 0, 0, 0, 0, 1, 1),
		(drawing, 738, 738, 0, 0, 0, 0, 1, 1),
		(drawing, 737, 737, 0, 0, 0, 0, 1, 1),
		(drawing, 736, 736, 0, 0, 0, 0, 1, 1),
		(drawing, 735, 735, 0, 0, 0, 0, 1, 1),
		(drawing, 734, 734, 0, 0, 0, 0, 1, 1),
		(drawing, 733, 733, 0, 0, 0, 0, 1, 1),
		(drawing, 732, 732, 0, 0, 0, 0, 1, 1),
		(drawing, 731, 731, 0, 0, 0, 0, 1, 1),
		(drawing, 730, 730, 0, 0, 0, 0, 1, 1),
		(drawing, 729, 729, 0, 0, 0, 0, 1, 1),
		(drawing, 728, 728, 0, 0, 0, 0, 1, 1),
		(drawing, 727, 727, 0, 0, 0, 0, 1, 1),
		(drawing, 726, 726, 0, 0, 0, 0, 1, 1),
		(drawing, 725, 725, 0, 0, 0, 0, 1, 1),
		(drawing, 724, 724, 0, 0, 0, 0, 1, 1),
		(drawing, 723, 723, 0, 0, 0, 0, 1, 1),
		(drawing, 722, 722, 0, 0, 0, 0, 1, 1),
		(drawing, 721, 721, 0, 0, 0, 0, 1, 1),
		(drawing, 720, 720, 0, 0, 0, 0, 1, 1),
		(drawing, 719, 719, 0, 0, 0, 0, 1, 1),
		(drawing, 718, 718, 0, 0, 0, 0, 1, 1),
		(drawing, 717, 717, 0, 0, 0, 0, 1, 1),
		(drawing, 716, 716, 0, 0, 0, 0, 1, 1),
		(drawing, 715, 715, 0, 0, 0, 0, 1, 1),
		(drawing, 714, 714, 0, 0, 0, 0, 1, 1),
		(drawing, 713, 713, 0, 0, 0, 0, 1, 1),
		(drawing, 712, 712, 0, 0, 0, 0, 1, 1),
		(drawing, 711, 711, 0, 0, 0, 0, 1, 1),
		(drawing, 710, 710, 0, 0, 0, 0, 1, 1),
		(drawing, 709, 709, 0, 0, 0, 0, 1, 1),
		(drawing, 708, 708, 0, 0, 0, 0, 1, 1),
		(drawing, 707, 707, 0, 0, 0, 0, 1, 1),
		(drawing, 706, 706, 0, 0, 0, 0, 1, 1),
		(drawing, 705, 705, 0, 0, 0, 0, 1, 1),
		(drawing, 704, 704, 0, 0, 0, 0, 1, 1),
		(drawing, 703, 703, 0, 0, 0, 0, 1, 1),
		(drawing, 702, 702, 0, 0, 0, 0, 1, 1),
		(drawing, 701, 701, 0, 0, 0, 0, 1, 1),
		(drawing, 700, 700, 0, 0, 0, 0, 1, 1),
		(drawing, 699, 699, 0, 0, 0, 0, 1, 1),
		(drawing, 698, 698, 0, 0, 0, 0, 1, 1),
		(drawing, 697, 697, 0, 0, 0, 0, 1, 1),
		(drawing, 696, 696, 0, 0, 0, 0, 1, 1),
		(drawing, 695, 695, 0, 0, 0, 0, 1, 1),
		(drawing, 694, 694, 0, 0, 0, 0, 1, 1),
		(drawing, 693, 693, 0, 0, 0, 0, 1, 1),
		(drawing, 692, 692, 0, 0, 0, 0, 1, 1),
		(drawing, 691, 691, 0, 0, 0, 0, 1, 1),
		(drawing, 690, 690, 0, 0, 0, 0, 1, 1),
		(drawing, 689, 689, 0, 0, 0, 0, 1, 1),
		(drawing, 688, 688, 0, 0, 0, 0, 1, 1),
		(drawing, 687, 687, 0, 0, 0, 0, 1, 1),
		(drawing, 686, 686, 0, 0, 0, 0, 1, 1),
		(drawing, 685, 685, 0, 0, 0, 0, 1, 1),
		(drawing, 684, 684, 0, 0, 0, 0, 1, 1),
		(drawing, 683, 683, 0, 0, 0, 0, 1, 1),
		(drawing, 682, 682, 0, 0, 0, 0, 1, 1),
		(drawing, 681, 681, 0, 0, 0, 0, 1, 1),
		(drawing, 680, 680, 0, 0, 0, 0, 1, 1),
		(drawing, 679, 679, 0, 0, 0, 0, 1, 1),
		(drawing, 678, 678, 0, 0, 0, 0, 1, 1),
		(drawing, 677, 677, 0, 0, 0, 0, 1, 1),
		(drawing, 676, 676, 0, 0, 0, 0, 1, 1),
		(drawing, 675, 675, 0, 0, 0, 0, 1, 1),
		(drawing, 674, 674, 0, 0, 0, 0, 1, 1),
		(drawing, 673, 673, 0, 0, 0, 0, 1, 1),
		(drawing, 672, 672, 0, 0, 0, 0, 1, 1),
		(drawing, 671, 671, 0, 0, 0, 0, 1, 1),
		(drawing, 670, 670, 0, 0, 0, 0, 1, 1),
		(drawing, 669, 669, 0, 0, 0, 0, 1, 1),
		(drawing, 668, 668, 0, 0, 0, 0, 1, 1),
		(drawing, 667, 667, 0, 0, 0, 0, 1, 1),
		(drawing, 666, 666, 0, 0, 0, 0, 1, 1),
		(drawing, 665, 665, 0, 0, 0, 0, 1, 1),
		(drawing, 664, 664, 0, 0, 0, 0, 1, 1),
		(drawing, 663, 663, 0, 0, 0, 0, 1, 1),
		(drawing, 662, 662, 0, 0, 0, 0, 1, 1),
		(drawing, 661, 661, 0, 0, 0, 0, 1, 1),
		(drawing, 660, 660, 0, 0, 0, 0, 1, 1),
		(drawing, 659, 659, 0, 0, 0, 0, 1, 1),
		(drawing, 658, 658, 0, 0, 0, 0, 1, 1),
		(drawing, 657, 657, 0, 0, 0, 0, 1, 1),
		(drawing, 656, 656, 0, 0, 0, 0, 1, 1),
		(drawing, 655, 655, 0, 0, 0, 0, 1, 1),
		(drawing, 654, 654, 0, 0, 0, 0, 1, 1),
		(drawing, 653, 653, 0, 0, 0, 0, 1, 1),
		(drawing, 652, 652, 0, 0, 0, 0, 1, 1),
		(drawing, 651, 651, 0, 0, 0, 0, 1, 1),
		(drawing, 650, 650, 0, 0, 0, 0, 1, 1),
		(drawing, 649, 649, 0, 0, 0, 0, 1, 1),
		(drawing, 648, 648, 0, 0, 0, 0, 1, 1),
		(drawing, 647, 647, 0, 0, 0, 0, 1, 1),
		(drawing, 646, 646, 0, 0, 0, 0, 1, 1),
		(drawing, 645, 645, 0, 0, 0, 0, 1, 1),
		(drawing, 644, 644, 0, 0, 0, 0, 1, 1),
		(drawing, 643, 643, 0, 0, 0, 0, 1, 1),
		(drawing, 642, 642, 0, 0, 0, 0, 1, 1),
		(drawing, 641, 641, 0, 0, 0, 0, 1, 1),
		(drawing, 640, 640, 0, 0, 0, 0, 1, 1),
		(drawing, 639, 639, 0, 0, 0, 0, 1, 1),
		(drawing, 638, 638, 0, 0, 0, 0, 1, 1),
		(drawing, 637, 637, 0, 0, 0, 0, 1, 1),
		(drawing, 636, 636, 0, 0, 0, 0, 1, 1),
		(drawing, 635, 635, 0, 0, 0, 0, 1, 1),
		(drawing, 634, 634, 0, 0, 0, 0, 1, 1),
		(drawing, 633, 633, 0, 0, 0, 0, 1, 1),
		(drawing, 632, 632, 0, 0, 0, 0, 1, 1),
		(drawing, 631, 631, 0, 0, 0, 0, 1, 1),
		(drawing, 630, 630, 0, 0, 0, 0, 1, 1),
		(drawing, 629, 629, 0, 0, 0, 0, 1, 1),
		(drawing, 628, 628, 0, 0, 0, 0, 1, 1),
		(drawing, 627, 627, 0, 0, 0, 0, 1, 1),
		(drawing, 626, 626, 0, 0, 0, 0, 1, 1),
		(drawing, 625, 625, 0, 0, 0, 0, 1, 1),
		(drawing, 624, 624, 0, 0, 0, 0, 1, 1),
		(drawing, 623, 623, 0, 0, 0, 0, 1, 1),
		(drawing, 622, 622, 0, 0, 0, 0, 1, 1),
		(drawing, 621, 621, 0, 0, 0, 0, 1, 1),
		(drawing, 620, 620, 0, 0, 0, 0, 1, 1),
		(drawing, 619, 619, 0, 0, 0, 0, 1, 1),
		(drawing, 618, 618, 0, 0, 0, 0, 1, 1),
		(drawing, 617, 617, 0, 0, 0, 0, 1, 1),
		(drawing, 616, 616, 0, 0, 0, 0, 1, 1),
		(drawing, 615, 615, 0, 0, 0, 0, 1, 1),
		(drawing, 614, 614, 0, 0, 0, 0, 1, 1),
		(drawing, 613, 613, 0, 0, 0, 0, 1, 1),
		(drawing, 612, 612, 0, 0, 0, 0, 1, 1),
		(drawing, 611, 611, 0, 0, 0, 0, 1, 1),
		(drawing, 610, 610, 0, 0, 0, 0, 1, 1),
		(drawing, 609, 609, 0, 0, 0, 0, 1, 1),
		(drawing, 608, 608, 0, 0, 0, 0, 1, 1),
		(drawing, 607, 607, 0, 0, 0, 0, 1, 1),
		(drawing, 606, 606, 0, 0, 0, 0, 1, 1),
		(drawing, 605, 605, 0, 0, 0, 0, 1, 1),
		(drawing, 604, 604, 0, 0, 0, 0, 1, 1),
		(drawing, 603, 603, 0, 0, 0, 0, 1, 1),
		(drawing, 602, 602, 0, 0, 0, 0, 1, 1),
		(drawing, 601, 601, 0, 0, 0, 0, 1, 1),
		(drawing, 600, 600, 0, 0, 0, 0, 1, 1),
		(drawing, 599, 599, 0, 0, 0, 0, 1, 1),
		(drawing, 598, 598, 0, 0, 0, 0, 1, 1),
		(drawing, 597, 597, 0, 0, 0, 0, 1, 1),
		(drawing, 596, 596, 0, 0, 0, 0, 1, 1),
		(drawing, 595, 595, 0, 0, 0, 0, 1, 1),
		(drawing, 594, 594, 0, 0, 0, 0, 1, 1),
		(drawing, 593, 593, 0, 0, 0, 0, 1, 1),
		(drawing, 592, 592, 0, 0, 0, 0, 1, 1),
		(drawing, 591, 591, 0, 0, 0, 0, 1, 1),
		(drawing, 590, 590, 0, 0, 0, 0, 1, 1),
		(drawing, 589, 589, 0, 0, 0, 0, 1, 1),
		(drawing, 588, 588, 0, 0, 0, 0, 1, 1),
		(drawing, 587, 587, 0, 0, 0, 0, 1, 1),
		(drawing, 586, 586, 0, 0, 0, 0, 1, 1),
		(drawing, 585, 585, 0, 0, 0, 0, 1, 1),
		(drawing, 584, 584, 0, 0, 0, 0, 1, 1),
		(drawing, 583, 583, 0, 0, 0, 0, 1, 1),
		(drawing, 582, 582, 0, 0, 0, 0, 1, 1),
		(drawing, 581, 581, 0, 0, 0, 0, 1, 1),
		(drawing, 580, 580, 0, 0, 0, 0, 1, 1),
		(drawing, 579, 579, 0, 0, 0, 0, 1, 1),
		(drawing, 578, 578, 0, 0, 0, 0, 1, 1),
		(drawing, 577, 577, 0, 0, 0, 0, 1, 1),
		(drawing, 576, 576, 0, 0, 0, 0, 1, 1),
		(drawing, 575, 575, 0, 0, 0, 0, 1, 1),
		(drawing, 574, 574, 0, 0, 0, 0, 1, 1),
		(drawing, 573, 573, 0, 0, 0, 0, 1, 1),
		(drawing, 572, 572, 0, 0, 0, 0, 1, 1),
		(drawing, 571, 571, 0, 0, 0, 0, 1, 1),
		(drawing, 570, 570, 0, 0, 0, 0, 1, 1),
		(drawing, 569, 569, 0, 0, 0, 0, 1, 1),
		(drawing, 568, 568, 0, 0, 0, 0, 1, 1),
		(drawing, 567, 567, 0, 0, 0, 0, 1, 1),
		(drawing, 566, 566, 0, 0, 0, 0, 1, 1),
		(drawing, 565, 565, 0, 0, 0, 0, 1, 1),
		(drawing, 564, 564, 0, 0, 0, 0, 1, 1),
		(drawing, 563, 563, 0, 0, 0, 0, 1, 1),
		(drawing, 562, 562, 0, 0, 0, 0, 1, 1),
		(drawing, 561, 561, 0, 0, 0, 0, 1, 1),
		(drawing, 560, 560, 0, 0, 0, 0, 1, 1),
		(drawing, 559, 559, 0, 0, 0, 0, 1, 1),
		(drawing, 558, 558, 0, 0, 0, 0, 1, 1),
		(drawing, 557, 557, 0, 0, 0, 0, 1, 1),
		(drawing, 556, 556, 0, 0, 0, 0, 1, 1),
		(drawing, 555, 555, 0, 0, 0, 0, 1, 1),
		(drawing, 554, 554, 0, 0, 0, 0, 1, 1),
		(drawing, 553, 553, 0, 0, 0, 0, 1, 1),
		(drawing, 552, 552, 0, 0, 0, 0, 1, 1),
		(drawing, 551, 551, 0, 0, 0, 0, 1, 1),
		(drawing, 550, 550, 0, 0, 0, 0, 1, 1),
		(drawing, 549, 549, 0, 0, 0, 0, 1, 1),
		(drawing, 548, 548, 0, 0, 0, 0, 1, 1),
		(drawing, 547, 547, 0, 0, 0, 0, 1, 1),
		(drawing, 546, 546, 0, 0, 0, 0, 1, 1),
		(drawing, 545, 545, 0, 0, 0, 0, 1, 1),
		(drawing, 544, 544, 0, 0, 0, 0, 1, 1),
		(drawing, 543, 543, 0, 0, 0, 0, 1, 1),
		(drawing, 542, 542, 0, 0, 0, 0, 1, 1),
		(drawing, 541, 541, 0, 0, 0, 0, 1, 1),
		(drawing, 540, 540, 0, 0, 0, 0, 1, 1),
		(drawing, 539, 539, 0, 0, 0, 0, 1, 1),
		(drawing, 538, 538, 0, 0, 0, 0, 1, 1),
		(drawing, 537, 537, 0, 0, 0, 0, 1, 1),
		(drawing, 536, 536, 0, 0, 0, 0, 1, 1),
		(drawing, 535, 535, 0, 0, 0, 0, 1, 1),
		(drawing, 534, 534, 0, 0, 0, 0, 1, 1),
		(drawing, 533, 533, 0, 0, 0, 0, 1, 1),
		(drawing, 532, 532, 0, 0, 0, 0, 1, 1),
		(drawing, 531, 531, 0, 0, 0, 0, 1, 1),
		(drawing, 530, 530, 0, 0, 0, 0, 1, 1),
		(drawing, 529, 529, 0, 0, 0, 0, 1, 1),
		(drawing, 528, 528, 0, 0, 0, 0, 1, 1),
		(drawing, 527, 527, 0, 0, 0, 0, 1, 1),
		(drawing, 526, 526, 0, 0, 0, 0, 1, 1),
		(drawing, 525, 525, 0, 0, 0, 0, 1, 1),
		(drawing, 524, 524, 0, 0, 0, 0, 1, 1),
		(drawing, 523, 523, 0, 0, 0, 0, 1, 1),
		(drawing, 522, 522, 0, 0, 0, 0, 1, 1),
		(drawing, 521, 521, 0, 0, 0, 0, 1, 1),
		(drawing, 520, 520, 0, 0, 0, 0, 1, 1),
		(drawing, 519, 519, 0, 0, 0, 0, 1, 1),
		(drawing, 518, 518, 0, 0, 0, 0, 1, 1),
		(drawing, 517, 517, 0, 0, 0, 0, 1, 1),
		(drawing, 516, 516, 0, 0, 0, 0, 1, 1),
		(drawing, 515, 515, 0, 0, 0, 0, 1, 1),
		(drawing, 514, 514, 0, 0, 0, 0, 1, 1),
		(drawing, 513, 513, 0, 0, 0, 0, 1, 1),
		(drawing, 512, 512, 0, 0, 0, 0, 1, 1),
		(drawing, 511, 511, 0, 0, 0, 0, 1, 1),
		(drawing, 510, 510, 0, 0, 0, 0, 1, 1),
		(drawing, 509, 509, 0, 0, 0, 0, 1, 1),
		(drawing, 508, 508, 0, 0, 0, 0, 1, 1),
		(drawing, 507, 507, 0, 0, 0, 0, 1, 1),
		(drawing, 506, 506, 0, 0, 0, 0, 1, 1),
		(drawing, 505, 505, 0, 0, 0, 0, 1, 1),
		(drawing, 504, 504, 0, 0, 0, 0, 1, 1),
		(drawing, 503, 503, 0, 0, 0, 0, 1, 1),
		(drawing, 502, 502, 0, 0, 0, 0, 1, 1),
		(drawing, 501, 501, 0, 0, 0, 0, 1, 1),
		(drawing, 500, 500, 0, 0, 0, 0, 1, 1),
		(drawing, 499, 499, 0, 0, 0, 0, 1, 1),
		(drawing, 498, 498, 0, 0, 0, 0, 1, 1),
		(drawing, 497, 497, 0, 0, 0, 0, 1, 1),
		(drawing, 496, 496, 0, 0, 0, 0, 1, 1),
		(drawing, 495, 495, 0, 0, 0, 0, 1, 1),
		(drawing, 494, 494, 0, 0, 0, 0, 1, 1),
		(drawing, 493, 493, 0, 0, 0, 0, 1, 1),
		(drawing, 492, 492, 0, 0, 0, 0, 1, 1),
		(drawing, 491, 491, 0, 0, 0, 0, 1, 1),
		(drawing, 490, 490, 0, 0, 0, 0, 1, 1),
		(drawing, 489, 489, 0, 0, 0, 0, 1, 1),
		(drawing, 488, 488, 0, 0, 0, 0, 1, 1),
		(drawing, 487, 487, 0, 0, 0, 0, 1, 1),
		(drawing, 486, 486, 0, 0, 0, 0, 1, 1),
		(drawing, 485, 485, 0, 0, 0, 0, 1, 1),
		(drawing, 484, 484, 0, 0, 0, 0, 1, 1),
		(drawing, 483, 483, 0, 0, 0, 0, 1, 1),
		(drawing, 482, 482, 0, 0, 0, 0, 1, 1),
		(drawing, 481, 481, 0, 0, 0, 0, 1, 1),
		(drawing, 480, 480, 0, 0, 0, 0, 1, 1),
		(drawing, 479, 479, 0, 0, 0, 0, 1, 1),
		(drawing, 478, 478, 0, 0, 0, 0, 1, 1),
		(drawing, 477, 477, 0, 0, 0, 0, 1, 1),
		(drawing, 476, 476, 0, 0, 0, 0, 1, 1),
		(drawing, 475, 475, 0, 0, 0, 0, 1, 1),
		(drawing, 474, 474, 0, 0, 0, 0, 1, 1),
		(drawing, 473, 473, 0, 0, 0, 0, 1, 1),
		(drawing, 472, 472, 0, 0, 0, 0, 1, 1),
		(drawing, 471, 471, 0, 0, 0, 0, 1, 1),
		(drawing, 470, 470, 0, 0, 0, 0, 1, 1),
		(drawing, 469, 469, 0, 0, 0, 0, 1, 1),
		(drawing, 468, 468, 0, 0, 0, 0, 1, 1),
		(drawing, 467, 467, 0, 0, 0, 0, 1, 1),
		(drawing, 466, 466, 0, 0, 0, 0, 1, 1),
		(drawing, 465, 465, 0, 0, 0, 0, 1, 1),
		(drawing, 464, 464, 0, 0, 0, 0, 1, 1),
		(drawing, 463, 463, 0, 0, 0, 0, 1, 1),
		(drawing, 462, 462, 0, 0, 0, 0, 1, 1),
		(drawing, 461, 461, 0, 0, 0, 0, 1, 1),
		(drawing, 460, 460, 0, 0, 0, 0, 1, 1),
		(drawing, 459, 459, 0, 0, 0, 0, 1, 1),
		(drawing, 458, 458, 0, 0, 0, 0, 1, 1),
		(drawing, 457, 457, 0, 0, 0, 0, 1, 1),
		(drawing, 456, 456, 0, 0, 0, 0, 1, 1),
		(drawing, 455, 455, 0, 0, 0, 0, 1, 1),
		(drawing, 454, 454, 0, 0, 0, 0, 1, 1),
		(drawing, 453, 453, 0, 0, 0, 0, 1, 1),
		(drawing, 452, 452, 0, 0, 0, 0, 1, 1),
		(drawing, 451, 451, 0, 0, 0, 0, 1, 1),
		(drawing, 450, 450, 0, 0, 0, 0, 1, 1),
		(drawing, 449, 449, 0, 0, 0, 0, 1, 1),
		(drawing, 448, 448, 0, 0, 0, 0, 1, 1),
		(drawing, 447, 447, 0, 0, 0, 0, 1, 1),
		(drawing, 446, 446, 0, 0, 0, 0, 1, 1),
		(drawing, 445, 445, 0, 0, 0, 0, 1, 1),
		(drawing, 444, 444, 0, 0, 0, 0, 1, 1),
		(drawing, 443, 443, 0, 0, 0, 0, 1, 1),
		(drawing, 442, 442, 0, 0, 0, 0, 1, 1),
		(drawing, 441, 441, 0, 0, 0, 0, 1, 1),
		(drawing, 440, 440, 0, 0, 0, 0, 1, 1),
		(drawing, 439, 439, 0, 0, 0, 0, 1, 1),
		(drawing, 438, 438, 0, 0, 0, 0, 1, 1),
		(drawing, 437, 437, 0, 0, 0, 0, 1, 1),
		(drawing, 436, 436, 0, 0, 0, 0, 1, 1),
		(drawing, 435, 435, 0, 0, 0, 0, 1, 1),
		(drawing, 434, 434, 0, 0, 0, 0, 1, 1),
		(drawing, 433, 433, 0, 0, 0, 0, 1, 1),
		(drawing, 432, 432, 0, 0, 0, 0, 1, 1),
		(drawing, 431, 431, 0, 0, 0, 0, 1, 1),
		(drawing, 430, 430, 0, 0, 0, 0, 1, 1),
		(drawing, 429, 429, 0, 0, 0, 0, 1, 1),
		(drawing, 428, 428, 0, 0, 0, 0, 1, 1),
		(drawing, 427, 427, 0, 0, 0, 0, 1, 1),
		(drawing, 426, 426, 0, 0, 0, 0, 1, 1),
		(drawing, 425, 425, 0, 0, 0, 0, 1, 1),
		(drawing, 424, 424, 0, 0, 0, 0, 1, 1),
		(drawing, 423, 423, 0, 0, 0, 0, 1, 1),
		(drawing, 422, 422, 0, 0, 0, 0, 1, 1),
		(drawing, 421, 421, 0, 0, 0, 0, 1, 1),
		(drawing, 420, 420, 0, 0, 0, 0, 1, 1),
		(drawing, 419, 419, 0, 0, 0, 0, 1, 1),
		(drawing, 418, 418, 0, 0, 0, 0, 1, 1),
		(drawing, 417, 417, 0, 0, 0, 0, 1, 1),
		(drawing, 416, 416, 0, 0, 0, 0, 1, 1),
		(drawing, 415, 415, 0, 0, 0, 0, 1, 1),
		(drawing, 414, 414, 0, 0, 0, 0, 1, 1),
		(drawing, 413, 413, 0, 0, 0, 0, 1, 1),
		(drawing, 412, 412, 0, 0, 0, 0, 1, 1),
		(drawing, 411, 411, 0, 0, 0, 0, 1, 1),
		(drawing, 410, 410, 0, 0, 0, 0, 1, 1),
		(drawing, 409, 409, 0, 0, 0, 0, 1, 1),
		(drawing, 408, 408, 0, 0, 0, 0, 1, 1),
		(drawing, 407, 407, 0, 0, 0, 0, 1, 1),
		(drawing, 406, 406, 0, 0, 0, 0, 1, 1),
		(drawing, 405, 405, 0, 0, 0, 0, 1, 1),
		(drawing, 404, 404, 0, 0, 0, 0, 1, 1),
		(drawing, 403, 403, 0, 0, 0, 0, 1, 1),
		(drawing, 402, 402, 0, 0, 0, 0, 1, 1),
		(drawing, 401, 401, 0, 0, 0, 0, 1, 1),
		(drawing, 400, 400, 0, 0, 0, 0, 1, 1),
		(drawing, 399, 399, 0, 0, 0, 0, 1, 1),
		(drawing, 398, 398, 0, 0, 0, 0, 1, 1),
		(drawing, 397, 397, 0, 0, 0, 0, 1, 1),
		(drawing, 396, 396, 0, 0, 0, 0, 1, 1),
		(drawing, 395, 395, 0, 0, 0, 0, 1, 1),
		(drawing, 394, 394, 0, 0, 0, 0, 1, 1),
		(drawing, 393, 393, 0, 0, 0, 0, 1, 1),
		(drawing, 392, 392, 0, 0, 0, 0, 1, 1),
		(drawing, 391, 391, 0, 0, 0, 0, 1, 1),
		(drawing, 390, 390, 0, 0, 0, 0, 1, 1),
		(drawing, 389, 389, 0, 0, 0, 0, 1, 1),
		(drawing, 388, 388, 0, 0, 0, 0, 1, 1),
		(drawing, 387, 387, 0, 0, 0, 0, 1, 1),
		(drawing, 386, 386, 0, 0, 0, 0, 1, 1),
		(drawing, 385, 385, 0, 0, 0, 0, 1, 1),
		(drawing, 384, 384, 0, 0, 0, 0, 1, 1),
		(drawing, 383, 383, 0, 0, 0, 0, 1, 1),
		(drawing, 382, 382, 0, 0, 0, 0, 1, 1),
		(drawing, 381, 381, 0, 0, 0, 0, 1, 1),
		(drawing, 380, 380, 0, 0, 0, 0, 1, 1),
		(drawing, 379, 379, 0, 0, 0, 0, 1, 1),
		(drawing, 378, 378, 0, 0, 0, 0, 1, 1),
		(drawing, 377, 377, 0, 0, 0, 0, 1, 1),
		(drawing, 376, 376, 0, 0, 0, 0, 1, 1),
		(drawing, 375, 375, 0, 0, 0, 0, 1, 1),
		(drawing, 374, 374, 0, 0, 0, 0, 1, 1),
		(drawing, 373, 373, 0, 0, 0, 0, 1, 1),
		(drawing, 372, 372, 0, 0, 0, 0, 1, 1),
		(drawing, 371, 371, 0, 0, 0, 0, 1, 1),
		(drawing, 370, 370, 0, 0, 0, 0, 1, 1),
		(drawing, 369, 369, 0, 0, 0, 0, 1, 1),
		(drawing, 368, 368, 0, 0, 0, 0, 1, 1),
		(drawing, 367, 367, 0, 0, 0, 0, 1, 1),
		(drawing, 366, 366, 0, 0, 0, 0, 1, 1),
		(drawing, 365, 365, 0, 0, 0, 0, 1, 1),
		(drawing, 364, 364, 0, 0, 0, 0, 1, 1),
		(drawing, 363, 363, 0, 0, 0, 0, 1, 1),
		(drawing, 362, 362, 0, 0, 0, 0, 1, 1),
		(drawing, 361, 361, 0, 0, 0, 0, 1, 1),
		(drawing, 360, 360, 0, 0, 0, 0, 1, 1),
		(drawing, 359, 359, 0, 0, 0, 0, 1, 1),
		(drawing, 358, 358, 0, 0, 0, 0, 1, 1),
		(drawing, 357, 357, 0, 0, 0, 0, 1, 1),
		(drawing, 356, 356, 0, 0, 0, 0, 1, 1),
		(drawing, 355, 355, 0, 0, 0, 0, 1, 1),
		(drawing, 354, 354, 0, 0, 0, 0, 1, 1),
		(drawing, 353, 353, 0, 0, 0, 0, 1, 1),
		(drawing, 352, 352, 0, 0, 0, 0, 1, 1),
		(drawing, 351, 351, 0, 0, 0, 0, 1, 1),
		(drawing, 350, 350, 0, 0, 0, 0, 1, 1),
		(drawing, 349, 349, 0, 0, 0, 0, 1, 1),
		(drawing, 348, 348, 0, 0, 0, 0, 1, 1),
		(drawing, 347, 347, 0, 0, 0, 0, 1, 1),
		(drawing, 346, 346, 0, 0, 0, 0, 1, 1),
		(drawing, 345, 345, 0, 0, 0, 0, 1, 1),
		(drawing, 344, 344, 0, 0, 0, 0, 1, 1),
		(drawing, 343, 343, 0, 0, 0, 0, 1, 1),
		(drawing, 342, 342, 0, 0, 0, 0, 1, 1),
		(drawing, 341, 341, 0, 0, 0, 0, 1, 1),
		(drawing, 340, 340, 0, 0, 0, 0, 1, 1),
		(drawing, 339, 339, 0, 0, 0, 0, 1, 1),
		(drawing, 338, 338, 0, 0, 0, 0, 1, 1),
		(drawing, 337, 337, 0, 0, 0, 0, 1, 1),
		(drawing, 336, 336, 0, 0, 0, 0, 1, 1),
		(drawing, 335, 335, 0, 0, 0, 0, 1, 1),
		(drawing, 334, 334, 0, 0, 0, 0, 1, 1),
		(drawing, 333, 333, 0, 0, 0, 0, 1, 1),
		(drawing, 332, 332, 0, 0, 0, 0, 1, 1),
		(drawing, 331, 331, 0, 0, 0, 0, 1, 1),
		(drawing, 330, 330, 0, 0, 0, 0, 1, 1),
		(drawing, 329, 329, 0, 0, 0, 0, 1, 1),
		(drawing, 328, 328, 0, 0, 0, 0, 1, 1),
		(drawing, 327, 327, 0, 0, 0, 0, 1, 1),
		(drawing, 326, 326, 0, 0, 0, 0, 1, 1),
		(drawing, 325, 325, 0, 0, 0, 0, 1, 1),
		(drawing, 324, 324, 0, 0, 0, 0, 1, 1),
		(drawing, 323, 323, 0, 0, 0, 0, 1, 1),
		(drawing, 322, 322, 0, 0, 0, 0, 1, 1),
		(drawing, 321, 321, 0, 0, 0, 0, 1, 1),
		(drawing, 320, 320, 0, 0, 0, 0, 1, 1),
		(drawing, 319, 319, 0, 0, 0, 0, 1, 1),
		(drawing, 318, 318, 0, 0, 0, 0, 1, 1),
		(drawing, 317, 317, 0, 0, 0, 0, 1, 1),
		(drawing, 316, 316, 0, 0, 0, 0, 1, 1),
		(drawing, 315, 315, 0, 0, 0, 0, 1, 1),
		(drawing, 314, 314, 0, 0, 0, 0, 1, 1),
		(drawing, 313, 313, 0, 0, 0, 0, 1, 1),
		(drawing, 312, 312, 0, 0, 0, 0, 1, 1),
		(drawing, 311, 311, 0, 0, 0, 0, 1, 1),
		(drawing, 310, 310, 0, 0, 0, 0, 1, 1),
		(drawing, 309, 309, 0, 0, 0, 0, 1, 1),
		(drawing, 308, 308, 0, 0, 0, 0, 1, 1),
		(drawing, 307, 307, 0, 0, 0, 0, 1, 1),
		(drawing, 306, 306, 0, 0, 0, 0, 1, 1),
		(drawing, 305, 305, 0, 0, 0, 0, 1, 1),
		(drawing, 304, 304, 0, 0, 0, 0, 1, 1),
		(drawing, 303, 303, 0, 0, 0, 0, 1, 1),
		(drawing, 302, 302, 0, 0, 0, 0, 1, 1),
		(drawing, 301, 301, 0, 0, 0, 0, 1, 1),
		(drawing, 300, 300, 0, 0, 0, 0, 1, 1),
		(drawing, 299, 299, 0, 0, 0, 0, 1, 1),
		(drawing, 298, 298, 0, 0, 0, 0, 1, 1),
		(drawing, 297, 297, 0, 0, 0, 0, 1, 1),
		(drawing, 296, 296, 0, 0, 0, 0, 1, 1),
		(drawing, 295, 295, 0, 0, 0, 0, 1, 1),
		(drawing, 294, 294, 0, 0, 0, 0, 1, 1),
		(drawing, 293, 293, 0, 0, 0, 0, 1, 1),
		(drawing, 292, 292, 0, 0, 0, 0, 1, 1),
		(drawing, 291, 291, 0, 0, 0, 0, 1, 1),
		(drawing, 290, 290, 0, 0, 0, 0, 1, 1),
		(drawing, 289, 289, 0, 0, 0, 0, 1, 1),
		(drawing, 288, 288, 0, 0, 0, 0, 1, 1),
		(drawing, 287, 287, 0, 0, 0, 0, 1, 1),
		(drawing, 286, 286, 0, 0, 0, 0, 1, 1),
		(drawing, 285, 285, 0, 0, 0, 0, 1, 1),
		(drawing, 284, 284, 0, 0, 0, 0, 1, 1),
		(drawing, 283, 283, 0, 0, 0, 0, 1, 1),
		(drawing, 282, 282, 0, 0, 0, 0, 1, 1),
		(drawing, 281, 281, 0, 0, 0, 0, 1, 1),
		(drawing, 280, 280, 0, 0, 0, 0, 1, 1),
		(drawing, 279, 279, 0, 0, 0, 0, 1, 1),
		(drawing, 278, 278, 0, 0, 0, 0, 1, 1),
		(drawing, 277, 277, 0, 0, 0, 0, 1, 1),
		(drawing, 276, 276, 0, 0, 0, 0, 1, 1),
		(drawing, 275, 275, 0, 0, 0, 0, 1, 1),
		(drawing, 274, 274, 0, 0, 0, 0, 1, 1),
		(drawing, 273, 273, 0, 0, 0, 0, 1, 1),
		(drawing, 272, 272, 0, 0, 0, 0, 1, 1),
		(drawing, 271, 271, 0, 0, 0, 0, 1, 1),
		(drawing, 270, 270, 0, 0, 0, 0, 1, 1),
		(drawing, 269, 269, 0, 0, 0, 0, 1, 1),
		(drawing, 268, 268, 0, 0, 0, 0, 1, 1),
		(drawing, 267, 267, 0, 0, 0, 0, 1, 1),
		(drawing, 266, 266, 0, 0, 0, 0, 1, 1),
		(drawing, 265, 265, 0, 0, 0, 0, 1, 1),
		(drawing, 264, 264, 0, 0, 0, 0, 1, 1),
		(drawing, 263, 263, 0, 0, 0, 0, 1, 1),
		(drawing, 262, 262, 0, 0, 0, 0, 1, 1),
		(drawing, 261, 261, 0, 0, 0, 0, 1, 1),
		(drawing, 260, 260, 0, 0, 0, 0, 1, 1),
		(drawing, 259, 259, 0, 0, 0, 0, 1, 1),
		(drawing, 258, 258, 0, 0, 0, 0, 1, 1),
		(drawing, 257, 257, 0, 0, 0, 0, 1, 1),
		(drawing, 256, 256, 0, 0, 0, 0, 1, 1),
		(drawing, 255, 255, 0, 0, 0, 0, 1, 1),
		(drawing, 254, 254, 0, 0, 0, 0, 1, 1),
		(drawing, 253, 253, 0, 0, 0, 0, 1, 1),
		(drawing, 252, 252, 0, 0, 0, 0, 1, 1),
		(drawing, 251, 251, 0, 0, 0, 0, 1, 1),
		(drawing, 250, 250, 0, 0, 0, 0, 1, 1),
		(drawing, 249, 249, 0, 0, 0, 0, 1, 1),
		(drawing, 248, 248, 0, 0, 0, 0, 1, 1),
		(drawing, 247, 247, 0, 0, 0, 0, 1, 1),
		(drawing, 246, 246, 0, 0, 0, 0, 1, 1),
		(drawing, 245, 245, 0, 0, 0, 0, 1, 1),
		(drawing, 244, 244, 0, 0, 0, 0, 1, 1),
		(drawing, 243, 243, 0, 0, 0, 0, 1, 1),
		(drawing, 242, 242, 0, 0, 0, 0, 1, 1),
		(drawing, 241, 241, 0, 0, 0, 0, 1, 1),
		(drawing, 240, 240, 0, 0, 0, 0, 1, 1),
		(drawing, 239, 239, 0, 0, 0, 0, 1, 1),
		(drawing, 238, 238, 0, 0, 0, 0, 1, 1),
		(drawing, 237, 237, 0, 0, 0, 0, 1, 1),
		(drawing, 236, 236, 0, 0, 0, 0, 1, 1),
		(drawing, 235, 235, 0, 0, 0, 0, 1, 1),
		(drawing, 234, 234, 0, 0, 0, 0, 1, 1),
		(drawing, 233, 233, 0, 0, 0, 0, 1, 1),
		(drawing, 232, 232, 0, 0, 0, 0, 1, 1),
		(drawing, 231, 231, 0, 0, 0, 0, 1, 1),
		(drawing, 230, 230, 0, 0, 0, 0, 1, 1),
		(drawing, 229, 229, 0, 0, 0, 0, 1, 1),
		(drawing, 228, 228, 0, 0, 0, 0, 1, 1),
		(drawing, 227, 227, 0, 0, 0, 0, 1, 1),
		(drawing, 226, 226, 0, 0, 0, 0, 1, 1),
		(drawing, 225, 225, 0, 0, 0, 0, 1, 1),
		(drawing, 224, 224, 0, 0, 0, 0, 1, 1),
		(drawing, 223, 223, 0, 0, 0, 0, 1, 1),
		(drawing, 222, 222, 0, 0, 0, 0, 1, 1),
		(drawing, 221, 221, 0, 0, 0, 0, 1, 1),
		(drawing, 220, 220, 0, 0, 0, 0, 1, 1),
		(drawing, 219, 219, 0, 0, 0, 0, 1, 1),
		(drawing, 218, 218, 0, 0, 0, 0, 1, 1),
		(drawing, 217, 217, 0, 0, 0, 0, 1, 1),
		(drawing, 216, 216, 0, 0, 0, 0, 1, 1),
		(drawing, 215, 215, 0, 0, 0, 0, 1, 1),
		(drawing, 214, 214, 0, 0, 0, 0, 1, 1),
		(drawing, 213, 213, 0, 0, 0, 0, 1, 1),
		(drawing, 212, 212, 0, 0, 0, 0, 1, 1),
		(drawing, 211, 211, 0, 0, 0, 0, 1, 1),
		(drawing, 210, 210, 0, 0, 0, 0, 1, 1),
		(drawing, 209, 209, 0, 0, 0, 0, 1, 1),
		(drawing, 208, 208, 0, 0, 0, 0, 1, 1),
		(drawing, 207, 207, 0, 0, 0, 0, 1, 1),
		(drawing, 206, 206, 0, 0, 0, 0, 1, 1),
		(drawing, 205, 205, 0, 0, 0, 0, 1, 1),
		(drawing, 204, 204, 0, 0, 0, 0, 1, 1),
		(drawing, 203, 203, 0, 0, 0, 0, 1, 1),
		(drawing, 202, 202, 0, 0, 0, 0, 1, 1),
		(drawing, 201, 201, 0, 0, 0, 0, 1, 1),
		(drawing, 200, 200, 0, 0, 0, 0, 1, 1),
		(drawing, 199, 199, 0, 0, 0, 0, 1, 1),
		(drawing, 198, 198, 0, 0, 0, 0, 1, 1),
		(drawing, 197, 197, 0, 0, 0, 0, 1, 1),
		(drawing, 196, 196, 0, 0, 0, 0, 1, 1),
		(drawing, 195, 195, 0, 0, 0, 0, 1, 1),
		(drawing, 194, 194, 0, 0, 0, 0, 1, 1),
		(drawing, 193, 193, 0, 0, 0, 0, 1, 1),
		(drawing, 192, 192, 0, 0, 0, 0, 1, 1),
		(drawing, 191, 191, 0, 0, 0, 0, 1, 1),
		(drawing, 190, 190, 0, 0, 0, 0, 1, 1),
		(drawing, 189, 189, 0, 0, 0, 0, 1, 1),
		(drawing, 188, 188, 0, 0, 0, 0, 1, 1),
		(drawing, 187, 187, 0, 0, 0, 0, 1, 1),
		(drawing, 186, 186, 0, 0, 0, 0, 1, 1),
		(drawing, 185, 185, 0, 0, 0, 0, 1, 1),
		(drawing, 184, 184, 0, 0, 0, 0, 1, 1),
		(drawing, 183, 183, 0, 0, 0, 0, 1, 1),
		(drawing, 182, 182, 0, 0, 0, 0, 1, 1),
		(drawing, 181, 181, 0, 0, 0, 0, 1, 1),
		(drawing, 180, 180, 0, 0, 0, 0, 1, 1),
		(drawing, 179, 179, 0, 0, 0, 0, 1, 1),
		(drawing, 178, 178, 0, 0, 0, 0, 1, 1),
		(drawing, 177, 177, 0, 0, 0, 0, 1, 1),
		(drawing, 176, 176, 0, 0, 0, 0, 1, 1),
		(drawing, 175, 175, 0, 0, 0, 0, 1, 1),
		(drawing, 174, 174, 0, 0, 0, 0, 1, 1),
		(drawing, 173, 173, 0, 0, 0, 0, 1, 1),
		(drawing, 172, 172, 0, 0, 0, 0, 1, 1),
		(drawing, 171, 171, 0, 0, 0, 0, 1, 1),
		(drawing, 170, 170, 0, 0, 0, 0, 1, 1),
		(drawing, 169, 169, 0, 0, 0, 0, 1, 1),
		(drawing, 168, 168, 0, 0, 0, 0, 1, 1),
		(drawing, 167, 167, 0, 0, 0, 0, 1, 1),
		(drawing, 166, 166, 0, 0, 0, 0, 1, 1),
		(drawing, 165, 165, 0, 0, 0, 0, 1, 1),
		(drawing, 164, 164, 0, 0, 0, 0, 1, 1),
		(drawing, 163, 163, 0, 0, 0, 0, 1, 1),
		(drawing, 162, 162, 0, 0, 0, 0, 1, 1),
		(drawing, 161, 161, 0, 0, 0, 0, 1, 1),
		(drawing, 160, 160, 0, 0, 0, 0, 1, 1),
		(drawing, 159, 159, 0, 0, 0, 0, 1, 1),
		(drawing, 158, 158, 0, 0, 0, 0, 1, 1),
		(drawing, 157, 157, 0, 0, 0, 0, 1, 1),
		(drawing, 156, 156, 0, 0, 0, 0, 1, 1),
		(drawing, 155, 155, 0, 0, 0, 0, 1, 1),
		(drawing, 154, 154, 0, 0, 0, 0, 1, 1),
		(drawing, 153, 153, 0, 0, 0, 0, 1, 1),
		(drawing, 152, 152, 0, 0, 0, 0, 1, 1),
		(drawing, 151, 151, 0, 0, 0, 0, 1, 1),
		(drawing, 150, 150, 0, 0, 0, 0, 1, 1),
		(drawing, 149, 149, 0, 0, 0, 0, 1, 1),
		(drawing, 148, 148, 0, 0, 0, 0, 1, 1),
		(drawing, 147, 147, 0, 0, 0, 0, 1, 1),
		(drawing, 146, 146, 0, 0, 0, 0, 1, 1),
		(drawing, 145, 145, 0, 0, 0, 0, 1, 1),
		(drawing, 144, 144, 0, 0, 0, 0, 1, 1),
		(drawing, 143, 143, 0, 0, 0, 0, 1, 1),
		(drawing, 142, 142, 0, 0, 0, 0, 1, 1),
		(drawing, 141, 141, 0, 0, 0, 0, 1, 1),
		(drawing, 140, 140, 0, 0, 0, 0, 1, 1),
		(drawing, 139, 139, 0, 0, 0, 0, 1, 1),
		(drawing, 138, 138, 0, 0, 0, 0, 1, 1),
		(drawing, 137, 137, 0, 0, 0, 0, 1, 1),
		(drawing, 136, 136, 0, 0, 0, 0, 1, 1),
		(drawing, 135, 135, 0, 0, 0, 0, 1, 1),
		(drawing, 134, 134, 0, 0, 0, 0, 1, 1),
		(drawing, 133, 133, 0, 0, 0, 0, 1, 1),
		(drawing, 132, 132, 0, 0, 0, 0, 1, 1),
		(drawing, 131, 131, 0, 0, 0, 0, 1, 1),
		(drawing, 130, 130, 0, 0, 0, 0, 1, 1),
		(drawing, 129, 129, 0, 0, 0, 0, 1, 1),
		(drawing, 128, 128, 0, 0, 0, 0, 1, 1),
		(drawing, 127, 127, 0, 0, 0, 0, 1, 1),
		(drawing, 126, 126, 0, 0, 0, 0, 1, 1),
		(drawing, 125, 125, 0, 0, 0, 0, 1, 1),
		(drawing, 124, 124, 0, 0, 0, 0, 1, 1),
		(drawing, 123, 123, 0, 0, 0, 0, 1, 1),
		(drawing, 122, 122, 0, 0, 0, 0, 1, 1),
		(drawing, 121, 121, 0, 0, 0, 0, 1, 1),
		(drawing, 120, 120, 0, 0, 0, 0, 1, 1),
		(drawing, 119, 119, 0, 0, 0, 0, 1, 1),
		(drawing, 118, 118, 0, 0, 0, 0, 1, 1),
		(drawing, 117, 117, 0, 0, 0, 0, 1, 1),
		(drawing, 116, 116, 0, 0, 0, 0, 1, 1),
		(drawing, 115, 115, 0, 0, 0, 0, 1, 1),
		(drawing, 114, 114, 0, 0, 0, 0, 1, 1),
		(drawing, 113, 113, 0, 0, 0, 0, 1, 1),
		(drawing, 112, 112, 0, 0, 0, 0, 1, 1),
		(drawing, 111, 111, 0, 0, 0, 0, 1, 1),
		(drawing, 110, 110, 0, 0, 0, 0, 1, 1),
		(drawing, 109, 109, 0, 0, 0, 0, 1, 1),
		(drawing, 108, 108, 0, 0, 0, 0, 1, 1),
		(drawing, 107, 107, 0, 0, 0, 0, 1, 1),
		(drawing, 106, 106, 0, 0, 0, 0, 1, 1),
		(drawing, 105, 105, 0, 0, 0, 0, 1, 1),
		(drawing, 104, 104, 0, 0, 0, 0, 1, 1),
		(drawing, 103, 103, 0, 0, 0, 0, 1, 1),
		(drawing, 102, 102, 0, 0, 0, 0, 1, 1),
		(drawing, 101, 101, 0, 0, 0, 0, 1, 1),
		(drawing, 100, 100, 0, 0, 0, 0, 1, 1),
		(drawing, 99, 99, 0, 0, 0, 0, 1, 1),
		(drawing, 98, 98, 0, 0, 0, 0, 1, 1),
		(drawing, 97, 97, 0, 0, 0, 0, 1, 1),
		(drawing, 96, 96, 0, 0, 0, 0, 1, 1),
		(drawing, 95, 95, 0, 0, 0, 0, 1, 1),
		(drawing, 94, 94, 0, 0, 0, 0, 1, 1),
		(drawing, 93, 93, 0, 0, 0, 0, 1, 1),
		(drawing, 92, 92, 0, 0, 0, 0, 1, 1),
		(drawing, 91, 91, 0, 0, 0, 0, 1, 1),
		(drawing, 90, 90, 0, 0, 0, 0, 1, 1),
		(drawing, 89, 89, 0, 0, 0, 0, 1, 1),
		(drawing, 88, 88, 0, 0, 0, 0, 1, 1),
		(drawing, 87, 87, 0, 0, 0, 0, 1, 1),
		(drawing, 86, 86, 0, 0, 0, 0, 1, 1),
		(drawing, 85, 85, 0, 0, 0, 0, 1, 1),
		(drawing, 84, 84, 0, 0, 0, 0, 1, 1),
		(drawing, 83, 83, 0, 0, 0, 0, 1, 1),
		(drawing, 82, 82, 0, 0, 0, 0, 1, 1),
		(drawing, 81, 81, 0, 0, 0, 0, 1, 1),
		(drawing, 80, 80, 0, 0, 0, 0, 1, 1),
		(drawing, 79, 79, 0, 0, 0, 0, 1, 1),
		(drawing, 78, 78, 0, 0, 0, 0, 1, 1),
		(drawing, 77, 77, 0, 0, 0, 0, 1, 1),
		(drawing, 76, 76, 0, 0, 0, 0, 1, 1),
		(drawing, 75, 75, 0, 0, 0, 0, 1, 1),
		(drawing, 74, 74, 0, 0, 0, 0, 1, 1),
		(drawing, 73, 73, 0, 0, 0, 0, 1, 1),
		(drawing, 72, 72, 0, 0, 0, 0, 1, 1),
		(drawing, 71, 71, 0, 0, 0, 0, 1, 1),
		(drawing, 70, 70, 0, 0, 0, 0, 1, 1),
		(drawing, 69, 69, 0, 0, 0, 0, 1, 1),
		(drawing, 68, 68, 0, 0, 0, 0, 1, 1),
		(drawing, 67, 67, 0, 0, 0, 0, 1, 1),
		(drawing, 66, 66, 0, 0, 0, 0, 1, 1),
		(drawing, 65, 65, 0, 0, 0, 0, 1, 1),
		(drawing, 64, 64, 0, 0, 0, 0, 1, 1),
		(drawing, 63, 63, 0, 0, 0, 0, 1, 1),
		(drawing, 62, 62, 0, 0, 0, 0, 1, 1),
		(drawing, 61, 61, 0, 0, 0, 0, 1, 1),
		(drawing, 60, 60, 0, 0, 0, 0, 1, 1),
		(drawing, 59, 59, 0, 0, 0, 0, 1, 1),
		(drawing, 58, 58, 0, 0, 0, 0, 1, 1),
		(drawing, 57, 57, 0, 0, 0, 0, 1, 1),
		(drawing, 56, 56, 0, 0, 0, 0, 1, 1),
		(drawing, 55, 55, 0, 0, 0, 0, 1, 1),
		(drawing, 54, 54, 0, 0, 0, 0, 1, 1),
		(drawing, 53, 53, 0, 0, 0, 0, 1, 1),
		(drawing, 52, 52, 0, 0, 0, 0, 1, 1),
		(drawing, 51, 51, 0, 0, 0, 0, 1, 1),
		(drawing, 50, 50, 0, 0, 0, 0, 1, 1),
		(drawing, 49, 49, 0, 0, 0, 0, 1, 1),
		(drawing, 48, 48, 0, 0, 0, 0, 1, 1),
		(drawing, 47, 47, 0, 0, 0, 0, 1, 1),
		(drawing, 46, 46, 0, 0, 0, 0, 1, 1),
		(drawing, 45, 45, 0, 0, 0, 0, 1, 1),
		(drawing, 44, 44, 0, 0, 0, 0, 1, 1),
		(drawing, 43, 43, 0, 0, 0, 0, 1, 1),
		(drawing, 42, 42, 0, 0, 0, 0, 1, 1),
		(drawing, 41, 41, 0, 0, 0, 0, 1, 1),
		(drawing, 40, 40, 0, 0, 0, 0, 1, 1),
		(drawing, 39, 39, 0, 0, 0, 0, 1, 1),
		(drawing, 38, 38, 0, 0, 0, 0, 1, 1),
		(drawing, 37, 37, 0, 0, 0, 0, 1, 1),
		(drawing, 36, 36, 0, 0, 0, 0, 1, 1),
		(drawing, 35, 35, 0, 0, 0, 0, 1, 1),
		(drawing, 34, 34, 0, 0, 0, 0, 1, 1),
		(drawing, 33, 33, 0, 0, 0, 0, 1, 1),
		(drawing, 32, 32, 0, 0, 0, 0, 1, 1),
		(drawing, 31, 31, 0, 0, 0, 0, 1, 1),
		(drawing, 30, 30, 0, 0, 0, 0, 1, 1),
		(drawing, 29, 29, 0, 0, 0, 0, 1, 1),
		(drawing, 28, 28, 0, 0, 0, 0, 1, 1),
		(drawing, 27, 27, 0, 0, 0, 0, 1, 1),
		(drawing, 26, 26, 0, 0, 0, 0, 1, 1),
		(drawing, 25, 25, 0, 0, 0, 0, 1, 1),
		(drawing, 24, 24, 0, 0, 0, 0, 1, 1),
		(drawing, 23, 23, 0, 0, 0, 0, 1, 1),
		(drawing, 22, 22, 0, 0, 0, 0, 1, 1),
		(drawing, 21, 21, 0, 0, 0, 0, 1, 1),
		(drawing, 20, 20, 0, 0, 0, 0, 1, 1),
		(drawing, 19, 19, 0, 0, 0, 0, 1, 1),
		(drawing, 18, 18, 0, 0, 0, 0, 1, 1),
		(drawing, 17, 17, 0, 0, 0, 0, 1, 1),
		(drawing, 16, 16, 0, 0, 0, 0, 1, 1),
		(drawing, 15, 15, 0, 0, 0, 0, 1, 1),
		(drawing, 14, 14, 0, 0, 0, 0, 1, 1),
		(drawing, 13, 13, 0, 0, 0, 0, 1, 1),
		(drawing, 12, 12, 0, 0, 0, 0, 1, 1),
		(drawing, 11, 11, 0, 0, 0, 0, 1, 1),
		(drawing, 10, 10, 0, 0, 0, 0, 1, 1),
		(drawing, 9, 9, 0, 0, 0, 0, 1, 1),
		(drawing, 8, 8, 0, 0, 0, 0, 1, 1),
		(drawing, 7, 7, 0, 0, 0, 0, 1, 1),
		(drawing, 6, 6, 0, 0, 0, 0, 1, 1),
		(drawing, 5, 5, 0, 0, 0, 0, 1, 1),
		(drawing, 4, 4, 0, 0, 0, 0, 1, 1),
		(drawing, 3, 3, 0, 0, 0, 0, 1, 1),
		(drawing, 2, 2, 0, 0, 0, 0, 1, 1),
		(drawing, 1, 1, 0, 0, 0, 0, 1, 1),
		(done, 0, 0, 0, 0, 0, 0, 1, 1)
	);
END PACKAGE ex4_data_pak;
