-- advanced test 5
-- draw line from (0,0) to (2048,2048)
-- NOTE * xin,yin are 12bits logic vectors
--------* 2048 in decimal is b1000,0000,0000

PACKAGE ex1_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 0, 0, 0),
		(start, 0, 0, 2048, 2048, 0),
		(drawing, 0, 0, 2048, 2048, 0),
		(drawing, 1, 1, 2048, 2048, 0),
		(drawing, 2, 2, 2048, 2048, 0),
		(drawing, 3, 3, 2048, 2048, 0),
		(drawing, 4, 4, 2048, 2048, 0),
		(drawing, 5, 5, 2048, 2048, 0),
		(drawing, 6, 6, 2048, 2048, 0),
		(drawing, 7, 7, 2048, 2048, 0),
		(drawing, 8, 8, 2048, 2048, 0),
		(drawing, 9, 9, 2048, 2048, 0),
		(drawing, 10, 10, 2048, 2048, 0),
		(drawing, 11, 11, 2048, 2048, 0),
		(drawing, 12, 12, 2048, 2048, 0),
		(drawing, 13, 13, 2048, 2048, 0),
		(drawing, 14, 14, 2048, 2048, 0),
		(drawing, 15, 15, 2048, 2048, 0),
		(drawing, 16, 16, 2048, 2048, 0),
		(drawing, 17, 17, 2048, 2048, 0),
		(drawing, 18, 18, 2048, 2048, 0),
		(drawing, 19, 19, 2048, 2048, 0),
		(drawing, 20, 20, 2048, 2048, 0),
		(drawing, 21, 21, 2048, 2048, 0),
		(drawing, 22, 22, 2048, 2048, 0),
		(drawing, 23, 23, 2048, 2048, 0),
		(drawing, 24, 24, 2048, 2048, 0),
		(drawing, 25, 25, 2048, 2048, 0),
		(drawing, 26, 26, 2048, 2048, 0),
		(drawing, 27, 27, 2048, 2048, 0),
		(drawing, 28, 28, 2048, 2048, 0),
		(drawing, 29, 29, 2048, 2048, 0),
		(drawing, 30, 30, 2048, 2048, 0),
		(drawing, 31, 31, 2048, 2048, 0),
		(drawing, 32, 32, 2048, 2048, 0),
		(drawing, 33, 33, 2048, 2048, 0),
		(drawing, 34, 34, 2048, 2048, 0),
		(drawing, 35, 35, 2048, 2048, 0),
		(drawing, 36, 36, 2048, 2048, 0),
		(drawing, 37, 37, 2048, 2048, 0),
		(drawing, 38, 38, 2048, 2048, 0),
		(drawing, 39, 39, 2048, 2048, 0),
		(drawing, 40, 40, 2048, 2048, 0),
		(drawing, 41, 41, 2048, 2048, 0),
		(drawing, 42, 42, 2048, 2048, 0),
		(drawing, 43, 43, 2048, 2048, 0),
		(drawing, 44, 44, 2048, 2048, 0),
		(drawing, 45, 45, 2048, 2048, 0),
		(drawing, 46, 46, 2048, 2048, 0),
		(drawing, 47, 47, 2048, 2048, 0),
		(drawing, 48, 48, 2048, 2048, 0),
		(drawing, 49, 49, 2048, 2048, 0),
		(drawing, 50, 50, 2048, 2048, 0),
		(drawing, 51, 51, 2048, 2048, 0),
		(drawing, 52, 52, 2048, 2048, 0),
		(drawing, 53, 53, 2048, 2048, 0),
		(drawing, 54, 54, 2048, 2048, 0),
		(drawing, 55, 55, 2048, 2048, 0),
		(drawing, 56, 56, 2048, 2048, 0),
		(drawing, 57, 57, 2048, 2048, 0),
		(drawing, 58, 58, 2048, 2048, 0),
		(drawing, 59, 59, 2048, 2048, 0),
		(drawing, 60, 60, 2048, 2048, 0),
		(drawing, 61, 61, 2048, 2048, 0),
		(drawing, 62, 62, 2048, 2048, 0),
		(drawing, 63, 63, 2048, 2048, 0),
		(drawing, 64, 64, 2048, 2048, 0),
		(drawing, 65, 65, 2048, 2048, 0),
		(drawing, 66, 66, 2048, 2048, 0),
		(drawing, 67, 67, 2048, 2048, 0),
		(drawing, 68, 68, 2048, 2048, 0),
		(drawing, 69, 69, 2048, 2048, 0),
		(drawing, 70, 70, 2048, 2048, 0),
		(drawing, 71, 71, 2048, 2048, 0),
		(drawing, 72, 72, 2048, 2048, 0),
		(drawing, 73, 73, 2048, 2048, 0),
		(drawing, 74, 74, 2048, 2048, 0),
		(drawing, 75, 75, 2048, 2048, 0),
		(drawing, 76, 76, 2048, 2048, 0),
		(drawing, 77, 77, 2048, 2048, 0),
		(drawing, 78, 78, 2048, 2048, 0),
		(drawing, 79, 79, 2048, 2048, 0),
		(drawing, 80, 80, 2048, 2048, 0),
		(drawing, 81, 81, 2048, 2048, 0),
		(drawing, 82, 82, 2048, 2048, 0),
		(drawing, 83, 83, 2048, 2048, 0),
		(drawing, 84, 84, 2048, 2048, 0),
		(drawing, 85, 85, 2048, 2048, 0),
		(drawing, 86, 86, 2048, 2048, 0),
		(drawing, 87, 87, 2048, 2048, 0),
		(drawing, 88, 88, 2048, 2048, 0),
		(drawing, 89, 89, 2048, 2048, 0),
		(drawing, 90, 90, 2048, 2048, 0),
		(drawing, 91, 91, 2048, 2048, 0),
		(drawing, 92, 92, 2048, 2048, 0),
		(drawing, 93, 93, 2048, 2048, 0),
		(drawing, 94, 94, 2048, 2048, 0),
		(drawing, 95, 95, 2048, 2048, 0),
		(drawing, 96, 96, 2048, 2048, 0),
		(drawing, 97, 97, 2048, 2048, 0),
		(drawing, 98, 98, 2048, 2048, 0),
		(drawing, 99, 99, 2048, 2048, 0),
		(drawing, 100, 100, 2048, 2048, 0),
		(drawing, 101, 101, 2048, 2048, 0),
		(drawing, 102, 102, 2048, 2048, 0),
		(drawing, 103, 103, 2048, 2048, 0),
		(drawing, 104, 104, 2048, 2048, 0),
		(drawing, 105, 105, 2048, 2048, 0),
		(drawing, 106, 106, 2048, 2048, 0),
		(drawing, 107, 107, 2048, 2048, 0),
		(drawing, 108, 108, 2048, 2048, 0),
		(drawing, 109, 109, 2048, 2048, 0),
		(drawing, 110, 110, 2048, 2048, 0),
		(drawing, 111, 111, 2048, 2048, 0),
		(drawing, 112, 112, 2048, 2048, 0),
		(drawing, 113, 113, 2048, 2048, 0),
		(drawing, 114, 114, 2048, 2048, 0),
		(drawing, 115, 115, 2048, 2048, 0),
		(drawing, 116, 116, 2048, 2048, 0),
		(drawing, 117, 117, 2048, 2048, 0),
		(drawing, 118, 118, 2048, 2048, 0),
		(drawing, 119, 119, 2048, 2048, 0),
		(drawing, 120, 120, 2048, 2048, 0),
		(drawing, 121, 121, 2048, 2048, 0),
		(drawing, 122, 122, 2048, 2048, 0),
		(drawing, 123, 123, 2048, 2048, 0),
		(drawing, 124, 124, 2048, 2048, 0),
		(drawing, 125, 125, 2048, 2048, 0),
		(drawing, 126, 126, 2048, 2048, 0),
		(drawing, 127, 127, 2048, 2048, 0),
		(drawing, 128, 128, 2048, 2048, 0),
		(drawing, 129, 129, 2048, 2048, 0),
		(drawing, 130, 130, 2048, 2048, 0),
		(drawing, 131, 131, 2048, 2048, 0),
		(drawing, 132, 132, 2048, 2048, 0),
		(drawing, 133, 133, 2048, 2048, 0),
		(drawing, 134, 134, 2048, 2048, 0),
		(drawing, 135, 135, 2048, 2048, 0),
		(drawing, 136, 136, 2048, 2048, 0),
		(drawing, 137, 137, 2048, 2048, 0),
		(drawing, 138, 138, 2048, 2048, 0),
		(drawing, 139, 139, 2048, 2048, 0),
		(drawing, 140, 140, 2048, 2048, 0),
		(drawing, 141, 141, 2048, 2048, 0),
		(drawing, 142, 142, 2048, 2048, 0),
		(drawing, 143, 143, 2048, 2048, 0),
		(drawing, 144, 144, 2048, 2048, 0),
		(drawing, 145, 145, 2048, 2048, 0),
		(drawing, 146, 146, 2048, 2048, 0),
		(drawing, 147, 147, 2048, 2048, 0),
		(drawing, 148, 148, 2048, 2048, 0),
		(drawing, 149, 149, 2048, 2048, 0),
		(drawing, 150, 150, 2048, 2048, 0),
		(drawing, 151, 151, 2048, 2048, 0),
		(drawing, 152, 152, 2048, 2048, 0),
		(drawing, 153, 153, 2048, 2048, 0),
		(drawing, 154, 154, 2048, 2048, 0),
		(drawing, 155, 155, 2048, 2048, 0),
		(drawing, 156, 156, 2048, 2048, 0),
		(drawing, 157, 157, 2048, 2048, 0),
		(drawing, 158, 158, 2048, 2048, 0),
		(drawing, 159, 159, 2048, 2048, 0),
		(drawing, 160, 160, 2048, 2048, 0),
		(drawing, 161, 161, 2048, 2048, 0),
		(drawing, 162, 162, 2048, 2048, 0),
		(drawing, 163, 163, 2048, 2048, 0),
		(drawing, 164, 164, 2048, 2048, 0),
		(drawing, 165, 165, 2048, 2048, 0),
		(drawing, 166, 166, 2048, 2048, 0),
		(drawing, 167, 167, 2048, 2048, 0),
		(drawing, 168, 168, 2048, 2048, 0),
		(drawing, 169, 169, 2048, 2048, 0),
		(drawing, 170, 170, 2048, 2048, 0),
		(drawing, 171, 171, 2048, 2048, 0),
		(drawing, 172, 172, 2048, 2048, 0),
		(drawing, 173, 173, 2048, 2048, 0),
		(drawing, 174, 174, 2048, 2048, 0),
		(drawing, 175, 175, 2048, 2048, 0),
		(drawing, 176, 176, 2048, 2048, 0),
		(drawing, 177, 177, 2048, 2048, 0),
		(drawing, 178, 178, 2048, 2048, 0),
		(drawing, 179, 179, 2048, 2048, 0),
		(drawing, 180, 180, 2048, 2048, 0),
		(drawing, 181, 181, 2048, 2048, 0),
		(drawing, 182, 182, 2048, 2048, 0),
		(drawing, 183, 183, 2048, 2048, 0),
		(drawing, 184, 184, 2048, 2048, 0),
		(drawing, 185, 185, 2048, 2048, 0),
		(drawing, 186, 186, 2048, 2048, 0),
		(drawing, 187, 187, 2048, 2048, 0),
		(drawing, 188, 188, 2048, 2048, 0),
		(drawing, 189, 189, 2048, 2048, 0),
		(drawing, 190, 190, 2048, 2048, 0),
		(drawing, 191, 191, 2048, 2048, 0),
		(drawing, 192, 192, 2048, 2048, 0),
		(drawing, 193, 193, 2048, 2048, 0),
		(drawing, 194, 194, 2048, 2048, 0),
		(drawing, 195, 195, 2048, 2048, 0),
		(drawing, 196, 196, 2048, 2048, 0),
		(drawing, 197, 197, 2048, 2048, 0),
		(drawing, 198, 198, 2048, 2048, 0),
		(drawing, 199, 199, 2048, 2048, 0),
		(drawing, 200, 200, 2048, 2048, 0),
		(drawing, 201, 201, 2048, 2048, 0),
		(drawing, 202, 202, 2048, 2048, 0),
		(drawing, 203, 203, 2048, 2048, 0),
		(drawing, 204, 204, 2048, 2048, 0),
		(drawing, 205, 205, 2048, 2048, 0),
		(drawing, 206, 206, 2048, 2048, 0),
		(drawing, 207, 207, 2048, 2048, 0),
		(drawing, 208, 208, 2048, 2048, 0),
		(drawing, 209, 209, 2048, 2048, 0),
		(drawing, 210, 210, 2048, 2048, 0),
		(drawing, 211, 211, 2048, 2048, 0),
		(drawing, 212, 212, 2048, 2048, 0),
		(drawing, 213, 213, 2048, 2048, 0),
		(drawing, 214, 214, 2048, 2048, 0),
		(drawing, 215, 215, 2048, 2048, 0),
		(drawing, 216, 216, 2048, 2048, 0),
		(drawing, 217, 217, 2048, 2048, 0),
		(drawing, 218, 218, 2048, 2048, 0),
		(drawing, 219, 219, 2048, 2048, 0),
		(drawing, 220, 220, 2048, 2048, 0),
		(drawing, 221, 221, 2048, 2048, 0),
		(drawing, 222, 222, 2048, 2048, 0),
		(drawing, 223, 223, 2048, 2048, 0),
		(drawing, 224, 224, 2048, 2048, 0),
		(drawing, 225, 225, 2048, 2048, 0),
		(drawing, 226, 226, 2048, 2048, 0),
		(drawing, 227, 227, 2048, 2048, 0),
		(drawing, 228, 228, 2048, 2048, 0),
		(drawing, 229, 229, 2048, 2048, 0),
		(drawing, 230, 230, 2048, 2048, 0),
		(drawing, 231, 231, 2048, 2048, 0),
		(drawing, 232, 232, 2048, 2048, 0),
		(drawing, 233, 233, 2048, 2048, 0),
		(drawing, 234, 234, 2048, 2048, 0),
		(drawing, 235, 235, 2048, 2048, 0),
		(drawing, 236, 236, 2048, 2048, 0),
		(drawing, 237, 237, 2048, 2048, 0),
		(drawing, 238, 238, 2048, 2048, 0),
		(drawing, 239, 239, 2048, 2048, 0),
		(drawing, 240, 240, 2048, 2048, 0),
		(drawing, 241, 241, 2048, 2048, 0),
		(drawing, 242, 242, 2048, 2048, 0),
		(drawing, 243, 243, 2048, 2048, 0),
		(drawing, 244, 244, 2048, 2048, 0),
		(drawing, 245, 245, 2048, 2048, 0),
		(drawing, 246, 246, 2048, 2048, 0),
		(drawing, 247, 247, 2048, 2048, 0),
		(drawing, 248, 248, 2048, 2048, 0),
		(drawing, 249, 249, 2048, 2048, 0),
		(drawing, 250, 250, 2048, 2048, 0),
		(drawing, 251, 251, 2048, 2048, 0),
		(drawing, 252, 252, 2048, 2048, 0),
		(drawing, 253, 253, 2048, 2048, 0),
		(drawing, 254, 254, 2048, 2048, 0),
		(drawing, 255, 255, 2048, 2048, 0),
		(drawing, 256, 256, 2048, 2048, 0),
		(drawing, 257, 257, 2048, 2048, 0),
		(drawing, 258, 258, 2048, 2048, 0),
		(drawing, 259, 259, 2048, 2048, 0),
		(drawing, 260, 260, 2048, 2048, 0),
		(drawing, 261, 261, 2048, 2048, 0),
		(drawing, 262, 262, 2048, 2048, 0),
		(drawing, 263, 263, 2048, 2048, 0),
		(drawing, 264, 264, 2048, 2048, 0),
		(drawing, 265, 265, 2048, 2048, 0),
		(drawing, 266, 266, 2048, 2048, 0),
		(drawing, 267, 267, 2048, 2048, 0),
		(drawing, 268, 268, 2048, 2048, 0),
		(drawing, 269, 269, 2048, 2048, 0),
		(drawing, 270, 270, 2048, 2048, 0),
		(drawing, 271, 271, 2048, 2048, 0),
		(drawing, 272, 272, 2048, 2048, 0),
		(drawing, 273, 273, 2048, 2048, 0),
		(drawing, 274, 274, 2048, 2048, 0),
		(drawing, 275, 275, 2048, 2048, 0),
		(drawing, 276, 276, 2048, 2048, 0),
		(drawing, 277, 277, 2048, 2048, 0),
		(drawing, 278, 278, 2048, 2048, 0),
		(drawing, 279, 279, 2048, 2048, 0),
		(drawing, 280, 280, 2048, 2048, 0),
		(drawing, 281, 281, 2048, 2048, 0),
		(drawing, 282, 282, 2048, 2048, 0),
		(drawing, 283, 283, 2048, 2048, 0),
		(drawing, 284, 284, 2048, 2048, 0),
		(drawing, 285, 285, 2048, 2048, 0),
		(drawing, 286, 286, 2048, 2048, 0),
		(drawing, 287, 287, 2048, 2048, 0),
		(drawing, 288, 288, 2048, 2048, 0),
		(drawing, 289, 289, 2048, 2048, 0),
		(drawing, 290, 290, 2048, 2048, 0),
		(drawing, 291, 291, 2048, 2048, 0),
		(drawing, 292, 292, 2048, 2048, 0),
		(drawing, 293, 293, 2048, 2048, 0),
		(drawing, 294, 294, 2048, 2048, 0),
		(drawing, 295, 295, 2048, 2048, 0),
		(drawing, 296, 296, 2048, 2048, 0),
		(drawing, 297, 297, 2048, 2048, 0),
		(drawing, 298, 298, 2048, 2048, 0),
		(drawing, 299, 299, 2048, 2048, 0),
		(drawing, 300, 300, 2048, 2048, 0),
		(drawing, 301, 301, 2048, 2048, 0),
		(drawing, 302, 302, 2048, 2048, 0),
		(drawing, 303, 303, 2048, 2048, 0),
		(drawing, 304, 304, 2048, 2048, 0),
		(drawing, 305, 305, 2048, 2048, 0),
		(drawing, 306, 306, 2048, 2048, 0),
		(drawing, 307, 307, 2048, 2048, 0),
		(drawing, 308, 308, 2048, 2048, 0),
		(drawing, 309, 309, 2048, 2048, 0),
		(drawing, 310, 310, 2048, 2048, 0),
		(drawing, 311, 311, 2048, 2048, 0),
		(drawing, 312, 312, 2048, 2048, 0),
		(drawing, 313, 313, 2048, 2048, 0),
		(drawing, 314, 314, 2048, 2048, 0),
		(drawing, 315, 315, 2048, 2048, 0),
		(drawing, 316, 316, 2048, 2048, 0),
		(drawing, 317, 317, 2048, 2048, 0),
		(drawing, 318, 318, 2048, 2048, 0),
		(drawing, 319, 319, 2048, 2048, 0),
		(drawing, 320, 320, 2048, 2048, 0),
		(drawing, 321, 321, 2048, 2048, 0),
		(drawing, 322, 322, 2048, 2048, 0),
		(drawing, 323, 323, 2048, 2048, 0),
		(drawing, 324, 324, 2048, 2048, 0),
		(drawing, 325, 325, 2048, 2048, 0),
		(drawing, 326, 326, 2048, 2048, 0),
		(drawing, 327, 327, 2048, 2048, 0),
		(drawing, 328, 328, 2048, 2048, 0),
		(drawing, 329, 329, 2048, 2048, 0),
		(drawing, 330, 330, 2048, 2048, 0),
		(drawing, 331, 331, 2048, 2048, 0),
		(drawing, 332, 332, 2048, 2048, 0),
		(drawing, 333, 333, 2048, 2048, 0),
		(drawing, 334, 334, 2048, 2048, 0),
		(drawing, 335, 335, 2048, 2048, 0),
		(drawing, 336, 336, 2048, 2048, 0),
		(drawing, 337, 337, 2048, 2048, 0),
		(drawing, 338, 338, 2048, 2048, 0),
		(drawing, 339, 339, 2048, 2048, 0),
		(drawing, 340, 340, 2048, 2048, 0),
		(drawing, 341, 341, 2048, 2048, 0),
		(drawing, 342, 342, 2048, 2048, 0),
		(drawing, 343, 343, 2048, 2048, 0),
		(drawing, 344, 344, 2048, 2048, 0),
		(drawing, 345, 345, 2048, 2048, 0),
		(drawing, 346, 346, 2048, 2048, 0),
		(drawing, 347, 347, 2048, 2048, 0),
		(drawing, 348, 348, 2048, 2048, 0),
		(drawing, 349, 349, 2048, 2048, 0),
		(drawing, 350, 350, 2048, 2048, 0),
		(drawing, 351, 351, 2048, 2048, 0),
		(drawing, 352, 352, 2048, 2048, 0),
		(drawing, 353, 353, 2048, 2048, 0),
		(drawing, 354, 354, 2048, 2048, 0),
		(drawing, 355, 355, 2048, 2048, 0),
		(drawing, 356, 356, 2048, 2048, 0),
		(drawing, 357, 357, 2048, 2048, 0),
		(drawing, 358, 358, 2048, 2048, 0),
		(drawing, 359, 359, 2048, 2048, 0),
		(drawing, 360, 360, 2048, 2048, 0),
		(drawing, 361, 361, 2048, 2048, 0),
		(drawing, 362, 362, 2048, 2048, 0),
		(drawing, 363, 363, 2048, 2048, 0),
		(drawing, 364, 364, 2048, 2048, 0),
		(drawing, 365, 365, 2048, 2048, 0),
		(drawing, 366, 366, 2048, 2048, 0),
		(drawing, 367, 367, 2048, 2048, 0),
		(drawing, 368, 368, 2048, 2048, 0),
		(drawing, 369, 369, 2048, 2048, 0),
		(drawing, 370, 370, 2048, 2048, 0),
		(drawing, 371, 371, 2048, 2048, 0),
		(drawing, 372, 372, 2048, 2048, 0),
		(drawing, 373, 373, 2048, 2048, 0),
		(drawing, 374, 374, 2048, 2048, 0),
		(drawing, 375, 375, 2048, 2048, 0),
		(drawing, 376, 376, 2048, 2048, 0),
		(drawing, 377, 377, 2048, 2048, 0),
		(drawing, 378, 378, 2048, 2048, 0),
		(drawing, 379, 379, 2048, 2048, 0),
		(drawing, 380, 380, 2048, 2048, 0),
		(drawing, 381, 381, 2048, 2048, 0),
		(drawing, 382, 382, 2048, 2048, 0),
		(drawing, 383, 383, 2048, 2048, 0),
		(drawing, 384, 384, 2048, 2048, 0),
		(drawing, 385, 385, 2048, 2048, 0),
		(drawing, 386, 386, 2048, 2048, 0),
		(drawing, 387, 387, 2048, 2048, 0),
		(drawing, 388, 388, 2048, 2048, 0),
		(drawing, 389, 389, 2048, 2048, 0),
		(drawing, 390, 390, 2048, 2048, 0),
		(drawing, 391, 391, 2048, 2048, 0),
		(drawing, 392, 392, 2048, 2048, 0),
		(drawing, 393, 393, 2048, 2048, 0),
		(drawing, 394, 394, 2048, 2048, 0),
		(drawing, 395, 395, 2048, 2048, 0),
		(drawing, 396, 396, 2048, 2048, 0),
		(drawing, 397, 397, 2048, 2048, 0),
		(drawing, 398, 398, 2048, 2048, 0),
		(drawing, 399, 399, 2048, 2048, 0),
		(drawing, 400, 400, 2048, 2048, 0),
		(drawing, 401, 401, 2048, 2048, 0),
		(drawing, 402, 402, 2048, 2048, 0),
		(drawing, 403, 403, 2048, 2048, 0),
		(drawing, 404, 404, 2048, 2048, 0),
		(drawing, 405, 405, 2048, 2048, 0),
		(drawing, 406, 406, 2048, 2048, 0),
		(drawing, 407, 407, 2048, 2048, 0),
		(drawing, 408, 408, 2048, 2048, 0),
		(drawing, 409, 409, 2048, 2048, 0),
		(drawing, 410, 410, 2048, 2048, 0),
		(drawing, 411, 411, 2048, 2048, 0),
		(drawing, 412, 412, 2048, 2048, 0),
		(drawing, 413, 413, 2048, 2048, 0),
		(drawing, 414, 414, 2048, 2048, 0),
		(drawing, 415, 415, 2048, 2048, 0),
		(drawing, 416, 416, 2048, 2048, 0),
		(drawing, 417, 417, 2048, 2048, 0),
		(drawing, 418, 418, 2048, 2048, 0),
		(drawing, 419, 419, 2048, 2048, 0),
		(drawing, 420, 420, 2048, 2048, 0),
		(drawing, 421, 421, 2048, 2048, 0),
		(drawing, 422, 422, 2048, 2048, 0),
		(drawing, 423, 423, 2048, 2048, 0),
		(drawing, 424, 424, 2048, 2048, 0),
		(drawing, 425, 425, 2048, 2048, 0),
		(drawing, 426, 426, 2048, 2048, 0),
		(drawing, 427, 427, 2048, 2048, 0),
		(drawing, 428, 428, 2048, 2048, 0),
		(drawing, 429, 429, 2048, 2048, 0),
		(drawing, 430, 430, 2048, 2048, 0),
		(drawing, 431, 431, 2048, 2048, 0),
		(drawing, 432, 432, 2048, 2048, 0),
		(drawing, 433, 433, 2048, 2048, 0),
		(drawing, 434, 434, 2048, 2048, 0),
		(drawing, 435, 435, 2048, 2048, 0),
		(drawing, 436, 436, 2048, 2048, 0),
		(drawing, 437, 437, 2048, 2048, 0),
		(drawing, 438, 438, 2048, 2048, 0),
		(drawing, 439, 439, 2048, 2048, 0),
		(drawing, 440, 440, 2048, 2048, 0),
		(drawing, 441, 441, 2048, 2048, 0),
		(drawing, 442, 442, 2048, 2048, 0),
		(drawing, 443, 443, 2048, 2048, 0),
		(drawing, 444, 444, 2048, 2048, 0),
		(drawing, 445, 445, 2048, 2048, 0),
		(drawing, 446, 446, 2048, 2048, 0),
		(drawing, 447, 447, 2048, 2048, 0),
		(drawing, 448, 448, 2048, 2048, 0),
		(drawing, 449, 449, 2048, 2048, 0),
		(drawing, 450, 450, 2048, 2048, 0),
		(drawing, 451, 451, 2048, 2048, 0),
		(drawing, 452, 452, 2048, 2048, 0),
		(drawing, 453, 453, 2048, 2048, 0),
		(drawing, 454, 454, 2048, 2048, 0),
		(drawing, 455, 455, 2048, 2048, 0),
		(drawing, 456, 456, 2048, 2048, 0),
		(drawing, 457, 457, 2048, 2048, 0),
		(drawing, 458, 458, 2048, 2048, 0),
		(drawing, 459, 459, 2048, 2048, 0),
		(drawing, 460, 460, 2048, 2048, 0),
		(drawing, 461, 461, 2048, 2048, 0),
		(drawing, 462, 462, 2048, 2048, 0),
		(drawing, 463, 463, 2048, 2048, 0),
		(drawing, 464, 464, 2048, 2048, 0),
		(drawing, 465, 465, 2048, 2048, 0),
		(drawing, 466, 466, 2048, 2048, 0),
		(drawing, 467, 467, 2048, 2048, 0),
		(drawing, 468, 468, 2048, 2048, 0),
		(drawing, 469, 469, 2048, 2048, 0),
		(drawing, 470, 470, 2048, 2048, 0),
		(drawing, 471, 471, 2048, 2048, 0),
		(drawing, 472, 472, 2048, 2048, 0),
		(drawing, 473, 473, 2048, 2048, 0),
		(drawing, 474, 474, 2048, 2048, 0),
		(drawing, 475, 475, 2048, 2048, 0),
		(drawing, 476, 476, 2048, 2048, 0),
		(drawing, 477, 477, 2048, 2048, 0),
		(drawing, 478, 478, 2048, 2048, 0),
		(drawing, 479, 479, 2048, 2048, 0),
		(drawing, 480, 480, 2048, 2048, 0),
		(drawing, 481, 481, 2048, 2048, 0),
		(drawing, 482, 482, 2048, 2048, 0),
		(drawing, 483, 483, 2048, 2048, 0),
		(drawing, 484, 484, 2048, 2048, 0),
		(drawing, 485, 485, 2048, 2048, 0),
		(drawing, 486, 486, 2048, 2048, 0),
		(drawing, 487, 487, 2048, 2048, 0),
		(drawing, 488, 488, 2048, 2048, 0),
		(drawing, 489, 489, 2048, 2048, 0),
		(drawing, 490, 490, 2048, 2048, 0),
		(drawing, 491, 491, 2048, 2048, 0),
		(drawing, 492, 492, 2048, 2048, 0),
		(drawing, 493, 493, 2048, 2048, 0),
		(drawing, 494, 494, 2048, 2048, 0),
		(drawing, 495, 495, 2048, 2048, 0),
		(drawing, 496, 496, 2048, 2048, 0),
		(drawing, 497, 497, 2048, 2048, 0),
		(drawing, 498, 498, 2048, 2048, 0),
		(drawing, 499, 499, 2048, 2048, 0),
		(drawing, 500, 500, 2048, 2048, 0),
		(drawing, 501, 501, 2048, 2048, 0),
		(drawing, 502, 502, 2048, 2048, 0),
		(drawing, 503, 503, 2048, 2048, 0),
		(drawing, 504, 504, 2048, 2048, 0),
		(drawing, 505, 505, 2048, 2048, 0),
		(drawing, 506, 506, 2048, 2048, 0),
		(drawing, 507, 507, 2048, 2048, 0),
		(drawing, 508, 508, 2048, 2048, 0),
		(drawing, 509, 509, 2048, 2048, 0),
		(drawing, 510, 510, 2048, 2048, 0),
		(drawing, 511, 511, 2048, 2048, 0),
		(drawing, 512, 512, 2048, 2048, 0),
		(drawing, 513, 513, 2048, 2048, 0),
		(drawing, 514, 514, 2048, 2048, 0),
		(drawing, 515, 515, 2048, 2048, 0),
		(drawing, 516, 516, 2048, 2048, 0),
		(drawing, 517, 517, 2048, 2048, 0),
		(drawing, 518, 518, 2048, 2048, 0),
		(drawing, 519, 519, 2048, 2048, 0),
		(drawing, 520, 520, 2048, 2048, 0),
		(drawing, 521, 521, 2048, 2048, 0),
		(drawing, 522, 522, 2048, 2048, 0),
		(drawing, 523, 523, 2048, 2048, 0),
		(drawing, 524, 524, 2048, 2048, 0),
		(drawing, 525, 525, 2048, 2048, 0),
		(drawing, 526, 526, 2048, 2048, 0),
		(drawing, 527, 527, 2048, 2048, 0),
		(drawing, 528, 528, 2048, 2048, 0),
		(drawing, 529, 529, 2048, 2048, 0),
		(drawing, 530, 530, 2048, 2048, 0),
		(drawing, 531, 531, 2048, 2048, 0),
		(drawing, 532, 532, 2048, 2048, 0),
		(drawing, 533, 533, 2048, 2048, 0),
		(drawing, 534, 534, 2048, 2048, 0),
		(drawing, 535, 535, 2048, 2048, 0),
		(drawing, 536, 536, 2048, 2048, 0),
		(drawing, 537, 537, 2048, 2048, 0),
		(drawing, 538, 538, 2048, 2048, 0),
		(drawing, 539, 539, 2048, 2048, 0),
		(drawing, 540, 540, 2048, 2048, 0),
		(drawing, 541, 541, 2048, 2048, 0),
		(drawing, 542, 542, 2048, 2048, 0),
		(drawing, 543, 543, 2048, 2048, 0),
		(drawing, 544, 544, 2048, 2048, 0),
		(drawing, 545, 545, 2048, 2048, 0),
		(drawing, 546, 546, 2048, 2048, 0),
		(drawing, 547, 547, 2048, 2048, 0),
		(drawing, 548, 548, 2048, 2048, 0),
		(drawing, 549, 549, 2048, 2048, 0),
		(drawing, 550, 550, 2048, 2048, 0),
		(drawing, 551, 551, 2048, 2048, 0),
		(drawing, 552, 552, 2048, 2048, 0),
		(drawing, 553, 553, 2048, 2048, 0),
		(drawing, 554, 554, 2048, 2048, 0),
		(drawing, 555, 555, 2048, 2048, 0),
		(drawing, 556, 556, 2048, 2048, 0),
		(drawing, 557, 557, 2048, 2048, 0),
		(drawing, 558, 558, 2048, 2048, 0),
		(drawing, 559, 559, 2048, 2048, 0),
		(drawing, 560, 560, 2048, 2048, 0),
		(drawing, 561, 561, 2048, 2048, 0),
		(drawing, 562, 562, 2048, 2048, 0),
		(drawing, 563, 563, 2048, 2048, 0),
		(drawing, 564, 564, 2048, 2048, 0),
		(drawing, 565, 565, 2048, 2048, 0),
		(drawing, 566, 566, 2048, 2048, 0),
		(drawing, 567, 567, 2048, 2048, 0),
		(drawing, 568, 568, 2048, 2048, 0),
		(drawing, 569, 569, 2048, 2048, 0),
		(drawing, 570, 570, 2048, 2048, 0),
		(drawing, 571, 571, 2048, 2048, 0),
		(drawing, 572, 572, 2048, 2048, 0),
		(drawing, 573, 573, 2048, 2048, 0),
		(drawing, 574, 574, 2048, 2048, 0),
		(drawing, 575, 575, 2048, 2048, 0),
		(drawing, 576, 576, 2048, 2048, 0),
		(drawing, 577, 577, 2048, 2048, 0),
		(drawing, 578, 578, 2048, 2048, 0),
		(drawing, 579, 579, 2048, 2048, 0),
		(drawing, 580, 580, 2048, 2048, 0),
		(drawing, 581, 581, 2048, 2048, 0),
		(drawing, 582, 582, 2048, 2048, 0),
		(drawing, 583, 583, 2048, 2048, 0),
		(drawing, 584, 584, 2048, 2048, 0),
		(drawing, 585, 585, 2048, 2048, 0),
		(drawing, 586, 586, 2048, 2048, 0),
		(drawing, 587, 587, 2048, 2048, 0),
		(drawing, 588, 588, 2048, 2048, 0),
		(drawing, 589, 589, 2048, 2048, 0),
		(drawing, 590, 590, 2048, 2048, 0),
		(drawing, 591, 591, 2048, 2048, 0),
		(drawing, 592, 592, 2048, 2048, 0),
		(drawing, 593, 593, 2048, 2048, 0),
		(drawing, 594, 594, 2048, 2048, 0),
		(drawing, 595, 595, 2048, 2048, 0),
		(drawing, 596, 596, 2048, 2048, 0),
		(drawing, 597, 597, 2048, 2048, 0),
		(drawing, 598, 598, 2048, 2048, 0),
		(drawing, 599, 599, 2048, 2048, 0),
		(drawing, 600, 600, 2048, 2048, 0),
		(drawing, 601, 601, 2048, 2048, 0),
		(drawing, 602, 602, 2048, 2048, 0),
		(drawing, 603, 603, 2048, 2048, 0),
		(drawing, 604, 604, 2048, 2048, 0),
		(drawing, 605, 605, 2048, 2048, 0),
		(drawing, 606, 606, 2048, 2048, 0),
		(drawing, 607, 607, 2048, 2048, 0),
		(drawing, 608, 608, 2048, 2048, 0),
		(drawing, 609, 609, 2048, 2048, 0),
		(drawing, 610, 610, 2048, 2048, 0),
		(drawing, 611, 611, 2048, 2048, 0),
		(drawing, 612, 612, 2048, 2048, 0),
		(drawing, 613, 613, 2048, 2048, 0),
		(drawing, 614, 614, 2048, 2048, 0),
		(drawing, 615, 615, 2048, 2048, 0),
		(drawing, 616, 616, 2048, 2048, 0),
		(drawing, 617, 617, 2048, 2048, 0),
		(drawing, 618, 618, 2048, 2048, 0),
		(drawing, 619, 619, 2048, 2048, 0),
		(drawing, 620, 620, 2048, 2048, 0),
		(drawing, 621, 621, 2048, 2048, 0),
		(drawing, 622, 622, 2048, 2048, 0),
		(drawing, 623, 623, 2048, 2048, 0),
		(drawing, 624, 624, 2048, 2048, 0),
		(drawing, 625, 625, 2048, 2048, 0),
		(drawing, 626, 626, 2048, 2048, 0),
		(drawing, 627, 627, 2048, 2048, 0),
		(drawing, 628, 628, 2048, 2048, 0),
		(drawing, 629, 629, 2048, 2048, 0),
		(drawing, 630, 630, 2048, 2048, 0),
		(drawing, 631, 631, 2048, 2048, 0),
		(drawing, 632, 632, 2048, 2048, 0),
		(drawing, 633, 633, 2048, 2048, 0),
		(drawing, 634, 634, 2048, 2048, 0),
		(drawing, 635, 635, 2048, 2048, 0),
		(drawing, 636, 636, 2048, 2048, 0),
		(drawing, 637, 637, 2048, 2048, 0),
		(drawing, 638, 638, 2048, 2048, 0),
		(drawing, 639, 639, 2048, 2048, 0),
		(drawing, 640, 640, 2048, 2048, 0),
		(drawing, 641, 641, 2048, 2048, 0),
		(drawing, 642, 642, 2048, 2048, 0),
		(drawing, 643, 643, 2048, 2048, 0),
		(drawing, 644, 644, 2048, 2048, 0),
		(drawing, 645, 645, 2048, 2048, 0),
		(drawing, 646, 646, 2048, 2048, 0),
		(drawing, 647, 647, 2048, 2048, 0),
		(drawing, 648, 648, 2048, 2048, 0),
		(drawing, 649, 649, 2048, 2048, 0),
		(drawing, 650, 650, 2048, 2048, 0),
		(drawing, 651, 651, 2048, 2048, 0),
		(drawing, 652, 652, 2048, 2048, 0),
		(drawing, 653, 653, 2048, 2048, 0),
		(drawing, 654, 654, 2048, 2048, 0),
		(drawing, 655, 655, 2048, 2048, 0),
		(drawing, 656, 656, 2048, 2048, 0),
		(drawing, 657, 657, 2048, 2048, 0),
		(drawing, 658, 658, 2048, 2048, 0),
		(drawing, 659, 659, 2048, 2048, 0),
		(drawing, 660, 660, 2048, 2048, 0),
		(drawing, 661, 661, 2048, 2048, 0),
		(drawing, 662, 662, 2048, 2048, 0),
		(drawing, 663, 663, 2048, 2048, 0),
		(drawing, 664, 664, 2048, 2048, 0),
		(drawing, 665, 665, 2048, 2048, 0),
		(drawing, 666, 666, 2048, 2048, 0),
		(drawing, 667, 667, 2048, 2048, 0),
		(drawing, 668, 668, 2048, 2048, 0),
		(drawing, 669, 669, 2048, 2048, 0),
		(drawing, 670, 670, 2048, 2048, 0),
		(drawing, 671, 671, 2048, 2048, 0),
		(drawing, 672, 672, 2048, 2048, 0),
		(drawing, 673, 673, 2048, 2048, 0),
		(drawing, 674, 674, 2048, 2048, 0),
		(drawing, 675, 675, 2048, 2048, 0),
		(drawing, 676, 676, 2048, 2048, 0),
		(drawing, 677, 677, 2048, 2048, 0),
		(drawing, 678, 678, 2048, 2048, 0),
		(drawing, 679, 679, 2048, 2048, 0),
		(drawing, 680, 680, 2048, 2048, 0),
		(drawing, 681, 681, 2048, 2048, 0),
		(drawing, 682, 682, 2048, 2048, 0),
		(drawing, 683, 683, 2048, 2048, 0),
		(drawing, 684, 684, 2048, 2048, 0),
		(drawing, 685, 685, 2048, 2048, 0),
		(drawing, 686, 686, 2048, 2048, 0),
		(drawing, 687, 687, 2048, 2048, 0),
		(drawing, 688, 688, 2048, 2048, 0),
		(drawing, 689, 689, 2048, 2048, 0),
		(drawing, 690, 690, 2048, 2048, 0),
		(drawing, 691, 691, 2048, 2048, 0),
		(drawing, 692, 692, 2048, 2048, 0),
		(drawing, 693, 693, 2048, 2048, 0),
		(drawing, 694, 694, 2048, 2048, 0),
		(drawing, 695, 695, 2048, 2048, 0),
		(drawing, 696, 696, 2048, 2048, 0),
		(drawing, 697, 697, 2048, 2048, 0),
		(drawing, 698, 698, 2048, 2048, 0),
		(drawing, 699, 699, 2048, 2048, 0),
		(drawing, 700, 700, 2048, 2048, 0),
		(drawing, 701, 701, 2048, 2048, 0),
		(drawing, 702, 702, 2048, 2048, 0),
		(drawing, 703, 703, 2048, 2048, 0),
		(drawing, 704, 704, 2048, 2048, 0),
		(drawing, 705, 705, 2048, 2048, 0),
		(drawing, 706, 706, 2048, 2048, 0),
		(drawing, 707, 707, 2048, 2048, 0),
		(drawing, 708, 708, 2048, 2048, 0),
		(drawing, 709, 709, 2048, 2048, 0),
		(drawing, 710, 710, 2048, 2048, 0),
		(drawing, 711, 711, 2048, 2048, 0),
		(drawing, 712, 712, 2048, 2048, 0),
		(drawing, 713, 713, 2048, 2048, 0),
		(drawing, 714, 714, 2048, 2048, 0),
		(drawing, 715, 715, 2048, 2048, 0),
		(drawing, 716, 716, 2048, 2048, 0),
		(drawing, 717, 717, 2048, 2048, 0),
		(drawing, 718, 718, 2048, 2048, 0),
		(drawing, 719, 719, 2048, 2048, 0),
		(drawing, 720, 720, 2048, 2048, 0),
		(drawing, 721, 721, 2048, 2048, 0),
		(drawing, 722, 722, 2048, 2048, 0),
		(drawing, 723, 723, 2048, 2048, 0),
		(drawing, 724, 724, 2048, 2048, 0),
		(drawing, 725, 725, 2048, 2048, 0),
		(drawing, 726, 726, 2048, 2048, 0),
		(drawing, 727, 727, 2048, 2048, 0),
		(drawing, 728, 728, 2048, 2048, 0),
		(drawing, 729, 729, 2048, 2048, 0),
		(drawing, 730, 730, 2048, 2048, 0),
		(drawing, 731, 731, 2048, 2048, 0),
		(drawing, 732, 732, 2048, 2048, 0),
		(drawing, 733, 733, 2048, 2048, 0),
		(drawing, 734, 734, 2048, 2048, 0),
		(drawing, 735, 735, 2048, 2048, 0),
		(drawing, 736, 736, 2048, 2048, 0),
		(drawing, 737, 737, 2048, 2048, 0),
		(drawing, 738, 738, 2048, 2048, 0),
		(drawing, 739, 739, 2048, 2048, 0),
		(drawing, 740, 740, 2048, 2048, 0),
		(drawing, 741, 741, 2048, 2048, 0),
		(drawing, 742, 742, 2048, 2048, 0),
		(drawing, 743, 743, 2048, 2048, 0),
		(drawing, 744, 744, 2048, 2048, 0),
		(drawing, 745, 745, 2048, 2048, 0),
		(drawing, 746, 746, 2048, 2048, 0),
		(drawing, 747, 747, 2048, 2048, 0),
		(drawing, 748, 748, 2048, 2048, 0),
		(drawing, 749, 749, 2048, 2048, 0),
		(drawing, 750, 750, 2048, 2048, 0),
		(drawing, 751, 751, 2048, 2048, 0),
		(drawing, 752, 752, 2048, 2048, 0),
		(drawing, 753, 753, 2048, 2048, 0),
		(drawing, 754, 754, 2048, 2048, 0),
		(drawing, 755, 755, 2048, 2048, 0),
		(drawing, 756, 756, 2048, 2048, 0),
		(drawing, 757, 757, 2048, 2048, 0),
		(drawing, 758, 758, 2048, 2048, 0),
		(drawing, 759, 759, 2048, 2048, 0),
		(drawing, 760, 760, 2048, 2048, 0),
		(drawing, 761, 761, 2048, 2048, 0),
		(drawing, 762, 762, 2048, 2048, 0),
		(drawing, 763, 763, 2048, 2048, 0),
		(drawing, 764, 764, 2048, 2048, 0),
		(drawing, 765, 765, 2048, 2048, 0),
		(drawing, 766, 766, 2048, 2048, 0),
		(drawing, 767, 767, 2048, 2048, 0),
		(drawing, 768, 768, 2048, 2048, 0),
		(drawing, 769, 769, 2048, 2048, 0),
		(drawing, 770, 770, 2048, 2048, 0),
		(drawing, 771, 771, 2048, 2048, 0),
		(drawing, 772, 772, 2048, 2048, 0),
		(drawing, 773, 773, 2048, 2048, 0),
		(drawing, 774, 774, 2048, 2048, 0),
		(drawing, 775, 775, 2048, 2048, 0),
		(drawing, 776, 776, 2048, 2048, 0),
		(drawing, 777, 777, 2048, 2048, 0),
		(drawing, 778, 778, 2048, 2048, 0),
		(drawing, 779, 779, 2048, 2048, 0),
		(drawing, 780, 780, 2048, 2048, 0),
		(drawing, 781, 781, 2048, 2048, 0),
		(drawing, 782, 782, 2048, 2048, 0),
		(drawing, 783, 783, 2048, 2048, 0),
		(drawing, 784, 784, 2048, 2048, 0),
		(drawing, 785, 785, 2048, 2048, 0),
		(drawing, 786, 786, 2048, 2048, 0),
		(drawing, 787, 787, 2048, 2048, 0),
		(drawing, 788, 788, 2048, 2048, 0),
		(drawing, 789, 789, 2048, 2048, 0),
		(drawing, 790, 790, 2048, 2048, 0),
		(drawing, 791, 791, 2048, 2048, 0),
		(drawing, 792, 792, 2048, 2048, 0),
		(drawing, 793, 793, 2048, 2048, 0),
		(drawing, 794, 794, 2048, 2048, 0),
		(drawing, 795, 795, 2048, 2048, 0),
		(drawing, 796, 796, 2048, 2048, 0),
		(drawing, 797, 797, 2048, 2048, 0),
		(drawing, 798, 798, 2048, 2048, 0),
		(drawing, 799, 799, 2048, 2048, 0),
		(drawing, 800, 800, 2048, 2048, 0),
		(drawing, 801, 801, 2048, 2048, 0),
		(drawing, 802, 802, 2048, 2048, 0),
		(drawing, 803, 803, 2048, 2048, 0),
		(drawing, 804, 804, 2048, 2048, 0),
		(drawing, 805, 805, 2048, 2048, 0),
		(drawing, 806, 806, 2048, 2048, 0),
		(drawing, 807, 807, 2048, 2048, 0),
		(drawing, 808, 808, 2048, 2048, 0),
		(drawing, 809, 809, 2048, 2048, 0),
		(drawing, 810, 810, 2048, 2048, 0),
		(drawing, 811, 811, 2048, 2048, 0),
		(drawing, 812, 812, 2048, 2048, 0),
		(drawing, 813, 813, 2048, 2048, 0),
		(drawing, 814, 814, 2048, 2048, 0),
		(drawing, 815, 815, 2048, 2048, 0),
		(drawing, 816, 816, 2048, 2048, 0),
		(drawing, 817, 817, 2048, 2048, 0),
		(drawing, 818, 818, 2048, 2048, 0),
		(drawing, 819, 819, 2048, 2048, 0),
		(drawing, 820, 820, 2048, 2048, 0),
		(drawing, 821, 821, 2048, 2048, 0),
		(drawing, 822, 822, 2048, 2048, 0),
		(drawing, 823, 823, 2048, 2048, 0),
		(drawing, 824, 824, 2048, 2048, 0),
		(drawing, 825, 825, 2048, 2048, 0),
		(drawing, 826, 826, 2048, 2048, 0),
		(drawing, 827, 827, 2048, 2048, 0),
		(drawing, 828, 828, 2048, 2048, 0),
		(drawing, 829, 829, 2048, 2048, 0),
		(drawing, 830, 830, 2048, 2048, 0),
		(drawing, 831, 831, 2048, 2048, 0),
		(drawing, 832, 832, 2048, 2048, 0),
		(drawing, 833, 833, 2048, 2048, 0),
		(drawing, 834, 834, 2048, 2048, 0),
		(drawing, 835, 835, 2048, 2048, 0),
		(drawing, 836, 836, 2048, 2048, 0),
		(drawing, 837, 837, 2048, 2048, 0),
		(drawing, 838, 838, 2048, 2048, 0),
		(drawing, 839, 839, 2048, 2048, 0),
		(drawing, 840, 840, 2048, 2048, 0),
		(drawing, 841, 841, 2048, 2048, 0),
		(drawing, 842, 842, 2048, 2048, 0),
		(drawing, 843, 843, 2048, 2048, 0),
		(drawing, 844, 844, 2048, 2048, 0),
		(drawing, 845, 845, 2048, 2048, 0),
		(drawing, 846, 846, 2048, 2048, 0),
		(drawing, 847, 847, 2048, 2048, 0),
		(drawing, 848, 848, 2048, 2048, 0),
		(drawing, 849, 849, 2048, 2048, 0),
		(drawing, 850, 850, 2048, 2048, 0),
		(drawing, 851, 851, 2048, 2048, 0),
		(drawing, 852, 852, 2048, 2048, 0),
		(drawing, 853, 853, 2048, 2048, 0),
		(drawing, 854, 854, 2048, 2048, 0),
		(drawing, 855, 855, 2048, 2048, 0),
		(drawing, 856, 856, 2048, 2048, 0),
		(drawing, 857, 857, 2048, 2048, 0),
		(drawing, 858, 858, 2048, 2048, 0),
		(drawing, 859, 859, 2048, 2048, 0),
		(drawing, 860, 860, 2048, 2048, 0),
		(drawing, 861, 861, 2048, 2048, 0),
		(drawing, 862, 862, 2048, 2048, 0),
		(drawing, 863, 863, 2048, 2048, 0),
		(drawing, 864, 864, 2048, 2048, 0),
		(drawing, 865, 865, 2048, 2048, 0),
		(drawing, 866, 866, 2048, 2048, 0),
		(drawing, 867, 867, 2048, 2048, 0),
		(drawing, 868, 868, 2048, 2048, 0),
		(drawing, 869, 869, 2048, 2048, 0),
		(drawing, 870, 870, 2048, 2048, 0),
		(drawing, 871, 871, 2048, 2048, 0),
		(drawing, 872, 872, 2048, 2048, 0),
		(drawing, 873, 873, 2048, 2048, 0),
		(drawing, 874, 874, 2048, 2048, 0),
		(drawing, 875, 875, 2048, 2048, 0),
		(drawing, 876, 876, 2048, 2048, 0),
		(drawing, 877, 877, 2048, 2048, 0),
		(drawing, 878, 878, 2048, 2048, 0),
		(drawing, 879, 879, 2048, 2048, 0),
		(drawing, 880, 880, 2048, 2048, 0),
		(drawing, 881, 881, 2048, 2048, 0),
		(drawing, 882, 882, 2048, 2048, 0),
		(drawing, 883, 883, 2048, 2048, 0),
		(drawing, 884, 884, 2048, 2048, 0),
		(drawing, 885, 885, 2048, 2048, 0),
		(drawing, 886, 886, 2048, 2048, 0),
		(drawing, 887, 887, 2048, 2048, 0),
		(drawing, 888, 888, 2048, 2048, 0),
		(drawing, 889, 889, 2048, 2048, 0),
		(drawing, 890, 890, 2048, 2048, 0),
		(drawing, 891, 891, 2048, 2048, 0),
		(drawing, 892, 892, 2048, 2048, 0),
		(drawing, 893, 893, 2048, 2048, 0),
		(drawing, 894, 894, 2048, 2048, 0),
		(drawing, 895, 895, 2048, 2048, 0),
		(drawing, 896, 896, 2048, 2048, 0),
		(drawing, 897, 897, 2048, 2048, 0),
		(drawing, 898, 898, 2048, 2048, 0),
		(drawing, 899, 899, 2048, 2048, 0),
		(drawing, 900, 900, 2048, 2048, 0),
		(drawing, 901, 901, 2048, 2048, 0),
		(drawing, 902, 902, 2048, 2048, 0),
		(drawing, 903, 903, 2048, 2048, 0),
		(drawing, 904, 904, 2048, 2048, 0),
		(drawing, 905, 905, 2048, 2048, 0),
		(drawing, 906, 906, 2048, 2048, 0),
		(drawing, 907, 907, 2048, 2048, 0),
		(drawing, 908, 908, 2048, 2048, 0),
		(drawing, 909, 909, 2048, 2048, 0),
		(drawing, 910, 910, 2048, 2048, 0),
		(drawing, 911, 911, 2048, 2048, 0),
		(drawing, 912, 912, 2048, 2048, 0),
		(drawing, 913, 913, 2048, 2048, 0),
		(drawing, 914, 914, 2048, 2048, 0),
		(drawing, 915, 915, 2048, 2048, 0),
		(drawing, 916, 916, 2048, 2048, 0),
		(drawing, 917, 917, 2048, 2048, 0),
		(drawing, 918, 918, 2048, 2048, 0),
		(drawing, 919, 919, 2048, 2048, 0),
		(drawing, 920, 920, 2048, 2048, 0),
		(drawing, 921, 921, 2048, 2048, 0),
		(drawing, 922, 922, 2048, 2048, 0),
		(drawing, 923, 923, 2048, 2048, 0),
		(drawing, 924, 924, 2048, 2048, 0),
		(drawing, 925, 925, 2048, 2048, 0),
		(drawing, 926, 926, 2048, 2048, 0),
		(drawing, 927, 927, 2048, 2048, 0),
		(drawing, 928, 928, 2048, 2048, 0),
		(drawing, 929, 929, 2048, 2048, 0),
		(drawing, 930, 930, 2048, 2048, 0),
		(drawing, 931, 931, 2048, 2048, 0),
		(drawing, 932, 932, 2048, 2048, 0),
		(drawing, 933, 933, 2048, 2048, 0),
		(drawing, 934, 934, 2048, 2048, 0),
		(drawing, 935, 935, 2048, 2048, 0),
		(drawing, 936, 936, 2048, 2048, 0),
		(drawing, 937, 937, 2048, 2048, 0),
		(drawing, 938, 938, 2048, 2048, 0),
		(drawing, 939, 939, 2048, 2048, 0),
		(drawing, 940, 940, 2048, 2048, 0),
		(drawing, 941, 941, 2048, 2048, 0),
		(drawing, 942, 942, 2048, 2048, 0),
		(drawing, 943, 943, 2048, 2048, 0),
		(drawing, 944, 944, 2048, 2048, 0),
		(drawing, 945, 945, 2048, 2048, 0),
		(drawing, 946, 946, 2048, 2048, 0),
		(drawing, 947, 947, 2048, 2048, 0),
		(drawing, 948, 948, 2048, 2048, 0),
		(drawing, 949, 949, 2048, 2048, 0),
		(drawing, 950, 950, 2048, 2048, 0),
		(drawing, 951, 951, 2048, 2048, 0),
		(drawing, 952, 952, 2048, 2048, 0),
		(drawing, 953, 953, 2048, 2048, 0),
		(drawing, 954, 954, 2048, 2048, 0),
		(drawing, 955, 955, 2048, 2048, 0),
		(drawing, 956, 956, 2048, 2048, 0),
		(drawing, 957, 957, 2048, 2048, 0),
		(drawing, 958, 958, 2048, 2048, 0),
		(drawing, 959, 959, 2048, 2048, 0),
		(drawing, 960, 960, 2048, 2048, 0),
		(drawing, 961, 961, 2048, 2048, 0),
		(drawing, 962, 962, 2048, 2048, 0),
		(drawing, 963, 963, 2048, 2048, 0),
		(drawing, 964, 964, 2048, 2048, 0),
		(drawing, 965, 965, 2048, 2048, 0),
		(drawing, 966, 966, 2048, 2048, 0),
		(drawing, 967, 967, 2048, 2048, 0),
		(drawing, 968, 968, 2048, 2048, 0),
		(drawing, 969, 969, 2048, 2048, 0),
		(drawing, 970, 970, 2048, 2048, 0),
		(drawing, 971, 971, 2048, 2048, 0),
		(drawing, 972, 972, 2048, 2048, 0),
		(drawing, 973, 973, 2048, 2048, 0),
		(drawing, 974, 974, 2048, 2048, 0),
		(drawing, 975, 975, 2048, 2048, 0),
		(drawing, 976, 976, 2048, 2048, 0),
		(drawing, 977, 977, 2048, 2048, 0),
		(drawing, 978, 978, 2048, 2048, 0),
		(drawing, 979, 979, 2048, 2048, 0),
		(drawing, 980, 980, 2048, 2048, 0),
		(drawing, 981, 981, 2048, 2048, 0),
		(drawing, 982, 982, 2048, 2048, 0),
		(drawing, 983, 983, 2048, 2048, 0),
		(drawing, 984, 984, 2048, 2048, 0),
		(drawing, 985, 985, 2048, 2048, 0),
		(drawing, 986, 986, 2048, 2048, 0),
		(drawing, 987, 987, 2048, 2048, 0),
		(drawing, 988, 988, 2048, 2048, 0),
		(drawing, 989, 989, 2048, 2048, 0),
		(drawing, 990, 990, 2048, 2048, 0),
		(drawing, 991, 991, 2048, 2048, 0),
		(drawing, 992, 992, 2048, 2048, 0),
		(drawing, 993, 993, 2048, 2048, 0),
		(drawing, 994, 994, 2048, 2048, 0),
		(drawing, 995, 995, 2048, 2048, 0),
		(drawing, 996, 996, 2048, 2048, 0),
		(drawing, 997, 997, 2048, 2048, 0),
		(drawing, 998, 998, 2048, 2048, 0),
		(drawing, 999, 999, 2048, 2048, 0),
		(drawing, 1000, 1000, 2048, 2048, 0),
		(drawing, 1001, 1001, 2048, 2048, 0),
		(drawing, 1002, 1002, 2048, 2048, 0),
		(drawing, 1003, 1003, 2048, 2048, 0),
		(drawing, 1004, 1004, 2048, 2048, 0),
		(drawing, 1005, 1005, 2048, 2048, 0),
		(drawing, 1006, 1006, 2048, 2048, 0),
		(drawing, 1007, 1007, 2048, 2048, 0),
		(drawing, 1008, 1008, 2048, 2048, 0),
		(drawing, 1009, 1009, 2048, 2048, 0),
		(drawing, 1010, 1010, 2048, 2048, 0),
		(drawing, 1011, 1011, 2048, 2048, 0),
		(drawing, 1012, 1012, 2048, 2048, 0),
		(drawing, 1013, 1013, 2048, 2048, 0),
		(drawing, 1014, 1014, 2048, 2048, 0),
		(drawing, 1015, 1015, 2048, 2048, 0),
		(drawing, 1016, 1016, 2048, 2048, 0),
		(drawing, 1017, 1017, 2048, 2048, 0),
		(drawing, 1018, 1018, 2048, 2048, 0),
		(drawing, 1019, 1019, 2048, 2048, 0),
		(drawing, 1020, 1020, 2048, 2048, 0),
		(drawing, 1021, 1021, 2048, 2048, 0),
		(drawing, 1022, 1022, 2048, 2048, 0),
		(drawing, 1023, 1023, 2048, 2048, 0),
		(drawing, 1024, 1024, 2048, 2048, 0),
		(drawing, 1025, 1025, 2048, 2048, 0),
		(drawing, 1026, 1026, 2048, 2048, 0),
		(drawing, 1027, 1027, 2048, 2048, 0),
		(drawing, 1028, 1028, 2048, 2048, 0),
		(drawing, 1029, 1029, 2048, 2048, 0),
		(drawing, 1030, 1030, 2048, 2048, 0),
		(drawing, 1031, 1031, 2048, 2048, 0),
		(drawing, 1032, 1032, 2048, 2048, 0),
		(drawing, 1033, 1033, 2048, 2048, 0),
		(drawing, 1034, 1034, 2048, 2048, 0),
		(drawing, 1035, 1035, 2048, 2048, 0),
		(drawing, 1036, 1036, 2048, 2048, 0),
		(drawing, 1037, 1037, 2048, 2048, 0),
		(drawing, 1038, 1038, 2048, 2048, 0),
		(drawing, 1039, 1039, 2048, 2048, 0),
		(drawing, 1040, 1040, 2048, 2048, 0),
		(drawing, 1041, 1041, 2048, 2048, 0),
		(drawing, 1042, 1042, 2048, 2048, 0),
		(drawing, 1043, 1043, 2048, 2048, 0),
		(drawing, 1044, 1044, 2048, 2048, 0),
		(drawing, 1045, 1045, 2048, 2048, 0),
		(drawing, 1046, 1046, 2048, 2048, 0),
		(drawing, 1047, 1047, 2048, 2048, 0),
		(drawing, 1048, 1048, 2048, 2048, 0),
		(drawing, 1049, 1049, 2048, 2048, 0),
		(drawing, 1050, 1050, 2048, 2048, 0),
		(drawing, 1051, 1051, 2048, 2048, 0),
		(drawing, 1052, 1052, 2048, 2048, 0),
		(drawing, 1053, 1053, 2048, 2048, 0),
		(drawing, 1054, 1054, 2048, 2048, 0),
		(drawing, 1055, 1055, 2048, 2048, 0),
		(drawing, 1056, 1056, 2048, 2048, 0),
		(drawing, 1057, 1057, 2048, 2048, 0),
		(drawing, 1058, 1058, 2048, 2048, 0),
		(drawing, 1059, 1059, 2048, 2048, 0),
		(drawing, 1060, 1060, 2048, 2048, 0),
		(drawing, 1061, 1061, 2048, 2048, 0),
		(drawing, 1062, 1062, 2048, 2048, 0),
		(drawing, 1063, 1063, 2048, 2048, 0),
		(drawing, 1064, 1064, 2048, 2048, 0),
		(drawing, 1065, 1065, 2048, 2048, 0),
		(drawing, 1066, 1066, 2048, 2048, 0),
		(drawing, 1067, 1067, 2048, 2048, 0),
		(drawing, 1068, 1068, 2048, 2048, 0),
		(drawing, 1069, 1069, 2048, 2048, 0),
		(drawing, 1070, 1070, 2048, 2048, 0),
		(drawing, 1071, 1071, 2048, 2048, 0),
		(drawing, 1072, 1072, 2048, 2048, 0),
		(drawing, 1073, 1073, 2048, 2048, 0),
		(drawing, 1074, 1074, 2048, 2048, 0),
		(drawing, 1075, 1075, 2048, 2048, 0),
		(drawing, 1076, 1076, 2048, 2048, 0),
		(drawing, 1077, 1077, 2048, 2048, 0),
		(drawing, 1078, 1078, 2048, 2048, 0),
		(drawing, 1079, 1079, 2048, 2048, 0),
		(drawing, 1080, 1080, 2048, 2048, 0),
		(drawing, 1081, 1081, 2048, 2048, 0),
		(drawing, 1082, 1082, 2048, 2048, 0),
		(drawing, 1083, 1083, 2048, 2048, 0),
		(drawing, 1084, 1084, 2048, 2048, 0),
		(drawing, 1085, 1085, 2048, 2048, 0),
		(drawing, 1086, 1086, 2048, 2048, 0),
		(drawing, 1087, 1087, 2048, 2048, 0),
		(drawing, 1088, 1088, 2048, 2048, 0),
		(drawing, 1089, 1089, 2048, 2048, 0),
		(drawing, 1090, 1090, 2048, 2048, 0),
		(drawing, 1091, 1091, 2048, 2048, 0),
		(drawing, 1092, 1092, 2048, 2048, 0),
		(drawing, 1093, 1093, 2048, 2048, 0),
		(drawing, 1094, 1094, 2048, 2048, 0),
		(drawing, 1095, 1095, 2048, 2048, 0),
		(drawing, 1096, 1096, 2048, 2048, 0),
		(drawing, 1097, 1097, 2048, 2048, 0),
		(drawing, 1098, 1098, 2048, 2048, 0),
		(drawing, 1099, 1099, 2048, 2048, 0),
		(drawing, 1100, 1100, 2048, 2048, 0),
		(drawing, 1101, 1101, 2048, 2048, 0),
		(drawing, 1102, 1102, 2048, 2048, 0),
		(drawing, 1103, 1103, 2048, 2048, 0),
		(drawing, 1104, 1104, 2048, 2048, 0),
		(drawing, 1105, 1105, 2048, 2048, 0),
		(drawing, 1106, 1106, 2048, 2048, 0),
		(drawing, 1107, 1107, 2048, 2048, 0),
		(drawing, 1108, 1108, 2048, 2048, 0),
		(drawing, 1109, 1109, 2048, 2048, 0),
		(drawing, 1110, 1110, 2048, 2048, 0),
		(drawing, 1111, 1111, 2048, 2048, 0),
		(drawing, 1112, 1112, 2048, 2048, 0),
		(drawing, 1113, 1113, 2048, 2048, 0),
		(drawing, 1114, 1114, 2048, 2048, 0),
		(drawing, 1115, 1115, 2048, 2048, 0),
		(drawing, 1116, 1116, 2048, 2048, 0),
		(drawing, 1117, 1117, 2048, 2048, 0),
		(drawing, 1118, 1118, 2048, 2048, 0),
		(drawing, 1119, 1119, 2048, 2048, 0),
		(drawing, 1120, 1120, 2048, 2048, 0),
		(drawing, 1121, 1121, 2048, 2048, 0),
		(drawing, 1122, 1122, 2048, 2048, 0),
		(drawing, 1123, 1123, 2048, 2048, 0),
		(drawing, 1124, 1124, 2048, 2048, 0),
		(drawing, 1125, 1125, 2048, 2048, 0),
		(drawing, 1126, 1126, 2048, 2048, 0),
		(drawing, 1127, 1127, 2048, 2048, 0),
		(drawing, 1128, 1128, 2048, 2048, 0),
		(drawing, 1129, 1129, 2048, 2048, 0),
		(drawing, 1130, 1130, 2048, 2048, 0),
		(drawing, 1131, 1131, 2048, 2048, 0),
		(drawing, 1132, 1132, 2048, 2048, 0),
		(drawing, 1133, 1133, 2048, 2048, 0),
		(drawing, 1134, 1134, 2048, 2048, 0),
		(drawing, 1135, 1135, 2048, 2048, 0),
		(drawing, 1136, 1136, 2048, 2048, 0),
		(drawing, 1137, 1137, 2048, 2048, 0),
		(drawing, 1138, 1138, 2048, 2048, 0),
		(drawing, 1139, 1139, 2048, 2048, 0),
		(drawing, 1140, 1140, 2048, 2048, 0),
		(drawing, 1141, 1141, 2048, 2048, 0),
		(drawing, 1142, 1142, 2048, 2048, 0),
		(drawing, 1143, 1143, 2048, 2048, 0),
		(drawing, 1144, 1144, 2048, 2048, 0),
		(drawing, 1145, 1145, 2048, 2048, 0),
		(drawing, 1146, 1146, 2048, 2048, 0),
		(drawing, 1147, 1147, 2048, 2048, 0),
		(drawing, 1148, 1148, 2048, 2048, 0),
		(drawing, 1149, 1149, 2048, 2048, 0),
		(drawing, 1150, 1150, 2048, 2048, 0),
		(drawing, 1151, 1151, 2048, 2048, 0),
		(drawing, 1152, 1152, 2048, 2048, 0),
		(drawing, 1153, 1153, 2048, 2048, 0),
		(drawing, 1154, 1154, 2048, 2048, 0),
		(drawing, 1155, 1155, 2048, 2048, 0),
		(drawing, 1156, 1156, 2048, 2048, 0),
		(drawing, 1157, 1157, 2048, 2048, 0),
		(drawing, 1158, 1158, 2048, 2048, 0),
		(drawing, 1159, 1159, 2048, 2048, 0),
		(drawing, 1160, 1160, 2048, 2048, 0),
		(drawing, 1161, 1161, 2048, 2048, 0),
		(drawing, 1162, 1162, 2048, 2048, 0),
		(drawing, 1163, 1163, 2048, 2048, 0),
		(drawing, 1164, 1164, 2048, 2048, 0),
		(drawing, 1165, 1165, 2048, 2048, 0),
		(drawing, 1166, 1166, 2048, 2048, 0),
		(drawing, 1167, 1167, 2048, 2048, 0),
		(drawing, 1168, 1168, 2048, 2048, 0),
		(drawing, 1169, 1169, 2048, 2048, 0),
		(drawing, 1170, 1170, 2048, 2048, 0),
		(drawing, 1171, 1171, 2048, 2048, 0),
		(drawing, 1172, 1172, 2048, 2048, 0),
		(drawing, 1173, 1173, 2048, 2048, 0),
		(drawing, 1174, 1174, 2048, 2048, 0),
		(drawing, 1175, 1175, 2048, 2048, 0),
		(drawing, 1176, 1176, 2048, 2048, 0),
		(drawing, 1177, 1177, 2048, 2048, 0),
		(drawing, 1178, 1178, 2048, 2048, 0),
		(drawing, 1179, 1179, 2048, 2048, 0),
		(drawing, 1180, 1180, 2048, 2048, 0),
		(drawing, 1181, 1181, 2048, 2048, 0),
		(drawing, 1182, 1182, 2048, 2048, 0),
		(drawing, 1183, 1183, 2048, 2048, 0),
		(drawing, 1184, 1184, 2048, 2048, 0),
		(drawing, 1185, 1185, 2048, 2048, 0),
		(drawing, 1186, 1186, 2048, 2048, 0),
		(drawing, 1187, 1187, 2048, 2048, 0),
		(drawing, 1188, 1188, 2048, 2048, 0),
		(drawing, 1189, 1189, 2048, 2048, 0),
		(drawing, 1190, 1190, 2048, 2048, 0),
		(drawing, 1191, 1191, 2048, 2048, 0),
		(drawing, 1192, 1192, 2048, 2048, 0),
		(drawing, 1193, 1193, 2048, 2048, 0),
		(drawing, 1194, 1194, 2048, 2048, 0),
		(drawing, 1195, 1195, 2048, 2048, 0),
		(drawing, 1196, 1196, 2048, 2048, 0),
		(drawing, 1197, 1197, 2048, 2048, 0),
		(drawing, 1198, 1198, 2048, 2048, 0),
		(drawing, 1199, 1199, 2048, 2048, 0),
		(drawing, 1200, 1200, 2048, 2048, 0),
		(drawing, 1201, 1201, 2048, 2048, 0),
		(drawing, 1202, 1202, 2048, 2048, 0),
		(drawing, 1203, 1203, 2048, 2048, 0),
		(drawing, 1204, 1204, 2048, 2048, 0),
		(drawing, 1205, 1205, 2048, 2048, 0),
		(drawing, 1206, 1206, 2048, 2048, 0),
		(drawing, 1207, 1207, 2048, 2048, 0),
		(drawing, 1208, 1208, 2048, 2048, 0),
		(drawing, 1209, 1209, 2048, 2048, 0),
		(drawing, 1210, 1210, 2048, 2048, 0),
		(drawing, 1211, 1211, 2048, 2048, 0),
		(drawing, 1212, 1212, 2048, 2048, 0),
		(drawing, 1213, 1213, 2048, 2048, 0),
		(drawing, 1214, 1214, 2048, 2048, 0),
		(drawing, 1215, 1215, 2048, 2048, 0),
		(drawing, 1216, 1216, 2048, 2048, 0),
		(drawing, 1217, 1217, 2048, 2048, 0),
		(drawing, 1218, 1218, 2048, 2048, 0),
		(drawing, 1219, 1219, 2048, 2048, 0),
		(drawing, 1220, 1220, 2048, 2048, 0),
		(drawing, 1221, 1221, 2048, 2048, 0),
		(drawing, 1222, 1222, 2048, 2048, 0),
		(drawing, 1223, 1223, 2048, 2048, 0),
		(drawing, 1224, 1224, 2048, 2048, 0),
		(drawing, 1225, 1225, 2048, 2048, 0),
		(drawing, 1226, 1226, 2048, 2048, 0),
		(drawing, 1227, 1227, 2048, 2048, 0),
		(drawing, 1228, 1228, 2048, 2048, 0),
		(drawing, 1229, 1229, 2048, 2048, 0),
		(drawing, 1230, 1230, 2048, 2048, 0),
		(drawing, 1231, 1231, 2048, 2048, 0),
		(drawing, 1232, 1232, 2048, 2048, 0),
		(drawing, 1233, 1233, 2048, 2048, 0),
		(drawing, 1234, 1234, 2048, 2048, 0),
		(drawing, 1235, 1235, 2048, 2048, 0),
		(drawing, 1236, 1236, 2048, 2048, 0),
		(drawing, 1237, 1237, 2048, 2048, 0),
		(drawing, 1238, 1238, 2048, 2048, 0),
		(drawing, 1239, 1239, 2048, 2048, 0),
		(drawing, 1240, 1240, 2048, 2048, 0),
		(drawing, 1241, 1241, 2048, 2048, 0),
		(drawing, 1242, 1242, 2048, 2048, 0),
		(drawing, 1243, 1243, 2048, 2048, 0),
		(drawing, 1244, 1244, 2048, 2048, 0),
		(drawing, 1245, 1245, 2048, 2048, 0),
		(drawing, 1246, 1246, 2048, 2048, 0),
		(drawing, 1247, 1247, 2048, 2048, 0),
		(drawing, 1248, 1248, 2048, 2048, 0),
		(drawing, 1249, 1249, 2048, 2048, 0),
		(drawing, 1250, 1250, 2048, 2048, 0),
		(drawing, 1251, 1251, 2048, 2048, 0),
		(drawing, 1252, 1252, 2048, 2048, 0),
		(drawing, 1253, 1253, 2048, 2048, 0),
		(drawing, 1254, 1254, 2048, 2048, 0),
		(drawing, 1255, 1255, 2048, 2048, 0),
		(drawing, 1256, 1256, 2048, 2048, 0),
		(drawing, 1257, 1257, 2048, 2048, 0),
		(drawing, 1258, 1258, 2048, 2048, 0),
		(drawing, 1259, 1259, 2048, 2048, 0),
		(drawing, 1260, 1260, 2048, 2048, 0),
		(drawing, 1261, 1261, 2048, 2048, 0),
		(drawing, 1262, 1262, 2048, 2048, 0),
		(drawing, 1263, 1263, 2048, 2048, 0),
		(drawing, 1264, 1264, 2048, 2048, 0),
		(drawing, 1265, 1265, 2048, 2048, 0),
		(drawing, 1266, 1266, 2048, 2048, 0),
		(drawing, 1267, 1267, 2048, 2048, 0),
		(drawing, 1268, 1268, 2048, 2048, 0),
		(drawing, 1269, 1269, 2048, 2048, 0),
		(drawing, 1270, 1270, 2048, 2048, 0),
		(drawing, 1271, 1271, 2048, 2048, 0),
		(drawing, 1272, 1272, 2048, 2048, 0),
		(drawing, 1273, 1273, 2048, 2048, 0),
		(drawing, 1274, 1274, 2048, 2048, 0),
		(drawing, 1275, 1275, 2048, 2048, 0),
		(drawing, 1276, 1276, 2048, 2048, 0),
		(drawing, 1277, 1277, 2048, 2048, 0),
		(drawing, 1278, 1278, 2048, 2048, 0),
		(drawing, 1279, 1279, 2048, 2048, 0),
		(drawing, 1280, 1280, 2048, 2048, 0),
		(drawing, 1281, 1281, 2048, 2048, 0),
		(drawing, 1282, 1282, 2048, 2048, 0),
		(drawing, 1283, 1283, 2048, 2048, 0),
		(drawing, 1284, 1284, 2048, 2048, 0),
		(drawing, 1285, 1285, 2048, 2048, 0),
		(drawing, 1286, 1286, 2048, 2048, 0),
		(drawing, 1287, 1287, 2048, 2048, 0),
		(drawing, 1288, 1288, 2048, 2048, 0),
		(drawing, 1289, 1289, 2048, 2048, 0),
		(drawing, 1290, 1290, 2048, 2048, 0),
		(drawing, 1291, 1291, 2048, 2048, 0),
		(drawing, 1292, 1292, 2048, 2048, 0),
		(drawing, 1293, 1293, 2048, 2048, 0),
		(drawing, 1294, 1294, 2048, 2048, 0),
		(drawing, 1295, 1295, 2048, 2048, 0),
		(drawing, 1296, 1296, 2048, 2048, 0),
		(drawing, 1297, 1297, 2048, 2048, 0),
		(drawing, 1298, 1298, 2048, 2048, 0),
		(drawing, 1299, 1299, 2048, 2048, 0),
		(drawing, 1300, 1300, 2048, 2048, 0),
		(drawing, 1301, 1301, 2048, 2048, 0),
		(drawing, 1302, 1302, 2048, 2048, 0),
		(drawing, 1303, 1303, 2048, 2048, 0),
		(drawing, 1304, 1304, 2048, 2048, 0),
		(drawing, 1305, 1305, 2048, 2048, 0),
		(drawing, 1306, 1306, 2048, 2048, 0),
		(drawing, 1307, 1307, 2048, 2048, 0),
		(drawing, 1308, 1308, 2048, 2048, 0),
		(drawing, 1309, 1309, 2048, 2048, 0),
		(drawing, 1310, 1310, 2048, 2048, 0),
		(drawing, 1311, 1311, 2048, 2048, 0),
		(drawing, 1312, 1312, 2048, 2048, 0),
		(drawing, 1313, 1313, 2048, 2048, 0),
		(drawing, 1314, 1314, 2048, 2048, 0),
		(drawing, 1315, 1315, 2048, 2048, 0),
		(drawing, 1316, 1316, 2048, 2048, 0),
		(drawing, 1317, 1317, 2048, 2048, 0),
		(drawing, 1318, 1318, 2048, 2048, 0),
		(drawing, 1319, 1319, 2048, 2048, 0),
		(drawing, 1320, 1320, 2048, 2048, 0),
		(drawing, 1321, 1321, 2048, 2048, 0),
		(drawing, 1322, 1322, 2048, 2048, 0),
		(drawing, 1323, 1323, 2048, 2048, 0),
		(drawing, 1324, 1324, 2048, 2048, 0),
		(drawing, 1325, 1325, 2048, 2048, 0),
		(drawing, 1326, 1326, 2048, 2048, 0),
		(drawing, 1327, 1327, 2048, 2048, 0),
		(drawing, 1328, 1328, 2048, 2048, 0),
		(drawing, 1329, 1329, 2048, 2048, 0),
		(drawing, 1330, 1330, 2048, 2048, 0),
		(drawing, 1331, 1331, 2048, 2048, 0),
		(drawing, 1332, 1332, 2048, 2048, 0),
		(drawing, 1333, 1333, 2048, 2048, 0),
		(drawing, 1334, 1334, 2048, 2048, 0),
		(drawing, 1335, 1335, 2048, 2048, 0),
		(drawing, 1336, 1336, 2048, 2048, 0),
		(drawing, 1337, 1337, 2048, 2048, 0),
		(drawing, 1338, 1338, 2048, 2048, 0),
		(drawing, 1339, 1339, 2048, 2048, 0),
		(drawing, 1340, 1340, 2048, 2048, 0),
		(drawing, 1341, 1341, 2048, 2048, 0),
		(drawing, 1342, 1342, 2048, 2048, 0),
		(drawing, 1343, 1343, 2048, 2048, 0),
		(drawing, 1344, 1344, 2048, 2048, 0),
		(drawing, 1345, 1345, 2048, 2048, 0),
		(drawing, 1346, 1346, 2048, 2048, 0),
		(drawing, 1347, 1347, 2048, 2048, 0),
		(drawing, 1348, 1348, 2048, 2048, 0),
		(drawing, 1349, 1349, 2048, 2048, 0),
		(drawing, 1350, 1350, 2048, 2048, 0),
		(drawing, 1351, 1351, 2048, 2048, 0),
		(drawing, 1352, 1352, 2048, 2048, 0),
		(drawing, 1353, 1353, 2048, 2048, 0),
		(drawing, 1354, 1354, 2048, 2048, 0),
		(drawing, 1355, 1355, 2048, 2048, 0),
		(drawing, 1356, 1356, 2048, 2048, 0),
		(drawing, 1357, 1357, 2048, 2048, 0),
		(drawing, 1358, 1358, 2048, 2048, 0),
		(drawing, 1359, 1359, 2048, 2048, 0),
		(drawing, 1360, 1360, 2048, 2048, 0),
		(drawing, 1361, 1361, 2048, 2048, 0),
		(drawing, 1362, 1362, 2048, 2048, 0),
		(drawing, 1363, 1363, 2048, 2048, 0),
		(drawing, 1364, 1364, 2048, 2048, 0),
		(drawing, 1365, 1365, 2048, 2048, 0),
		(drawing, 1366, 1366, 2048, 2048, 0),
		(drawing, 1367, 1367, 2048, 2048, 0),
		(drawing, 1368, 1368, 2048, 2048, 0),
		(drawing, 1369, 1369, 2048, 2048, 0),
		(drawing, 1370, 1370, 2048, 2048, 0),
		(drawing, 1371, 1371, 2048, 2048, 0),
		(drawing, 1372, 1372, 2048, 2048, 0),
		(drawing, 1373, 1373, 2048, 2048, 0),
		(drawing, 1374, 1374, 2048, 2048, 0),
		(drawing, 1375, 1375, 2048, 2048, 0),
		(drawing, 1376, 1376, 2048, 2048, 0),
		(drawing, 1377, 1377, 2048, 2048, 0),
		(drawing, 1378, 1378, 2048, 2048, 0),
		(drawing, 1379, 1379, 2048, 2048, 0),
		(drawing, 1380, 1380, 2048, 2048, 0),
		(drawing, 1381, 1381, 2048, 2048, 0),
		(drawing, 1382, 1382, 2048, 2048, 0),
		(drawing, 1383, 1383, 2048, 2048, 0),
		(drawing, 1384, 1384, 2048, 2048, 0),
		(drawing, 1385, 1385, 2048, 2048, 0),
		(drawing, 1386, 1386, 2048, 2048, 0),
		(drawing, 1387, 1387, 2048, 2048, 0),
		(drawing, 1388, 1388, 2048, 2048, 0),
		(drawing, 1389, 1389, 2048, 2048, 0),
		(drawing, 1390, 1390, 2048, 2048, 0),
		(drawing, 1391, 1391, 2048, 2048, 0),
		(drawing, 1392, 1392, 2048, 2048, 0),
		(drawing, 1393, 1393, 2048, 2048, 0),
		(drawing, 1394, 1394, 2048, 2048, 0),
		(drawing, 1395, 1395, 2048, 2048, 0),
		(drawing, 1396, 1396, 2048, 2048, 0),
		(drawing, 1397, 1397, 2048, 2048, 0),
		(drawing, 1398, 1398, 2048, 2048, 0),
		(drawing, 1399, 1399, 2048, 2048, 0),
		(drawing, 1400, 1400, 2048, 2048, 0),
		(drawing, 1401, 1401, 2048, 2048, 0),
		(drawing, 1402, 1402, 2048, 2048, 0),
		(drawing, 1403, 1403, 2048, 2048, 0),
		(drawing, 1404, 1404, 2048, 2048, 0),
		(drawing, 1405, 1405, 2048, 2048, 0),
		(drawing, 1406, 1406, 2048, 2048, 0),
		(drawing, 1407, 1407, 2048, 2048, 0),
		(drawing, 1408, 1408, 2048, 2048, 0),
		(drawing, 1409, 1409, 2048, 2048, 0),
		(drawing, 1410, 1410, 2048, 2048, 0),
		(drawing, 1411, 1411, 2048, 2048, 0),
		(drawing, 1412, 1412, 2048, 2048, 0),
		(drawing, 1413, 1413, 2048, 2048, 0),
		(drawing, 1414, 1414, 2048, 2048, 0),
		(drawing, 1415, 1415, 2048, 2048, 0),
		(drawing, 1416, 1416, 2048, 2048, 0),
		(drawing, 1417, 1417, 2048, 2048, 0),
		(drawing, 1418, 1418, 2048, 2048, 0),
		(drawing, 1419, 1419, 2048, 2048, 0),
		(drawing, 1420, 1420, 2048, 2048, 0),
		(drawing, 1421, 1421, 2048, 2048, 0),
		(drawing, 1422, 1422, 2048, 2048, 0),
		(drawing, 1423, 1423, 2048, 2048, 0),
		(drawing, 1424, 1424, 2048, 2048, 0),
		(drawing, 1425, 1425, 2048, 2048, 0),
		(drawing, 1426, 1426, 2048, 2048, 0),
		(drawing, 1427, 1427, 2048, 2048, 0),
		(drawing, 1428, 1428, 2048, 2048, 0),
		(drawing, 1429, 1429, 2048, 2048, 0),
		(drawing, 1430, 1430, 2048, 2048, 0),
		(drawing, 1431, 1431, 2048, 2048, 0),
		(drawing, 1432, 1432, 2048, 2048, 0),
		(drawing, 1433, 1433, 2048, 2048, 0),
		(drawing, 1434, 1434, 2048, 2048, 0),
		(drawing, 1435, 1435, 2048, 2048, 0),
		(drawing, 1436, 1436, 2048, 2048, 0),
		(drawing, 1437, 1437, 2048, 2048, 0),
		(drawing, 1438, 1438, 2048, 2048, 0),
		(drawing, 1439, 1439, 2048, 2048, 0),
		(drawing, 1440, 1440, 2048, 2048, 0),
		(drawing, 1441, 1441, 2048, 2048, 0),
		(drawing, 1442, 1442, 2048, 2048, 0),
		(drawing, 1443, 1443, 2048, 2048, 0),
		(drawing, 1444, 1444, 2048, 2048, 0),
		(drawing, 1445, 1445, 2048, 2048, 0),
		(drawing, 1446, 1446, 2048, 2048, 0),
		(drawing, 1447, 1447, 2048, 2048, 0),
		(drawing, 1448, 1448, 2048, 2048, 0),
		(drawing, 1449, 1449, 2048, 2048, 0),
		(drawing, 1450, 1450, 2048, 2048, 0),
		(drawing, 1451, 1451, 2048, 2048, 0),
		(drawing, 1452, 1452, 2048, 2048, 0),
		(drawing, 1453, 1453, 2048, 2048, 0),
		(drawing, 1454, 1454, 2048, 2048, 0),
		(drawing, 1455, 1455, 2048, 2048, 0),
		(drawing, 1456, 1456, 2048, 2048, 0),
		(drawing, 1457, 1457, 2048, 2048, 0),
		(drawing, 1458, 1458, 2048, 2048, 0),
		(drawing, 1459, 1459, 2048, 2048, 0),
		(drawing, 1460, 1460, 2048, 2048, 0),
		(drawing, 1461, 1461, 2048, 2048, 0),
		(drawing, 1462, 1462, 2048, 2048, 0),
		(drawing, 1463, 1463, 2048, 2048, 0),
		(drawing, 1464, 1464, 2048, 2048, 0),
		(drawing, 1465, 1465, 2048, 2048, 0),
		(drawing, 1466, 1466, 2048, 2048, 0),
		(drawing, 1467, 1467, 2048, 2048, 0),
		(drawing, 1468, 1468, 2048, 2048, 0),
		(drawing, 1469, 1469, 2048, 2048, 0),
		(drawing, 1470, 1470, 2048, 2048, 0),
		(drawing, 1471, 1471, 2048, 2048, 0),
		(drawing, 1472, 1472, 2048, 2048, 0),
		(drawing, 1473, 1473, 2048, 2048, 0),
		(drawing, 1474, 1474, 2048, 2048, 0),
		(drawing, 1475, 1475, 2048, 2048, 0),
		(drawing, 1476, 1476, 2048, 2048, 0),
		(drawing, 1477, 1477, 2048, 2048, 0),
		(drawing, 1478, 1478, 2048, 2048, 0),
		(drawing, 1479, 1479, 2048, 2048, 0),
		(drawing, 1480, 1480, 2048, 2048, 0),
		(drawing, 1481, 1481, 2048, 2048, 0),
		(drawing, 1482, 1482, 2048, 2048, 0),
		(drawing, 1483, 1483, 2048, 2048, 0),
		(drawing, 1484, 1484, 2048, 2048, 0),
		(drawing, 1485, 1485, 2048, 2048, 0),
		(drawing, 1486, 1486, 2048, 2048, 0),
		(drawing, 1487, 1487, 2048, 2048, 0),
		(drawing, 1488, 1488, 2048, 2048, 0),
		(drawing, 1489, 1489, 2048, 2048, 0),
		(drawing, 1490, 1490, 2048, 2048, 0),
		(drawing, 1491, 1491, 2048, 2048, 0),
		(drawing, 1492, 1492, 2048, 2048, 0),
		(drawing, 1493, 1493, 2048, 2048, 0),
		(drawing, 1494, 1494, 2048, 2048, 0),
		(drawing, 1495, 1495, 2048, 2048, 0),
		(drawing, 1496, 1496, 2048, 2048, 0),
		(drawing, 1497, 1497, 2048, 2048, 0),
		(drawing, 1498, 1498, 2048, 2048, 0),
		(drawing, 1499, 1499, 2048, 2048, 0),
		(drawing, 1500, 1500, 2048, 2048, 0),
		(drawing, 1501, 1501, 2048, 2048, 0),
		(drawing, 1502, 1502, 2048, 2048, 0),
		(drawing, 1503, 1503, 2048, 2048, 0),
		(drawing, 1504, 1504, 2048, 2048, 0),
		(drawing, 1505, 1505, 2048, 2048, 0),
		(drawing, 1506, 1506, 2048, 2048, 0),
		(drawing, 1507, 1507, 2048, 2048, 0),
		(drawing, 1508, 1508, 2048, 2048, 0),
		(drawing, 1509, 1509, 2048, 2048, 0),
		(drawing, 1510, 1510, 2048, 2048, 0),
		(drawing, 1511, 1511, 2048, 2048, 0),
		(drawing, 1512, 1512, 2048, 2048, 0),
		(drawing, 1513, 1513, 2048, 2048, 0),
		(drawing, 1514, 1514, 2048, 2048, 0),
		(drawing, 1515, 1515, 2048, 2048, 0),
		(drawing, 1516, 1516, 2048, 2048, 0),
		(drawing, 1517, 1517, 2048, 2048, 0),
		(drawing, 1518, 1518, 2048, 2048, 0),
		(drawing, 1519, 1519, 2048, 2048, 0),
		(drawing, 1520, 1520, 2048, 2048, 0),
		(drawing, 1521, 1521, 2048, 2048, 0),
		(drawing, 1522, 1522, 2048, 2048, 0),
		(drawing, 1523, 1523, 2048, 2048, 0),
		(drawing, 1524, 1524, 2048, 2048, 0),
		(drawing, 1525, 1525, 2048, 2048, 0),
		(drawing, 1526, 1526, 2048, 2048, 0),
		(drawing, 1527, 1527, 2048, 2048, 0),
		(drawing, 1528, 1528, 2048, 2048, 0),
		(drawing, 1529, 1529, 2048, 2048, 0),
		(drawing, 1530, 1530, 2048, 2048, 0),
		(drawing, 1531, 1531, 2048, 2048, 0),
		(drawing, 1532, 1532, 2048, 2048, 0),
		(drawing, 1533, 1533, 2048, 2048, 0),
		(drawing, 1534, 1534, 2048, 2048, 0),
		(drawing, 1535, 1535, 2048, 2048, 0),
		(drawing, 1536, 1536, 2048, 2048, 0),
		(drawing, 1537, 1537, 2048, 2048, 0),
		(drawing, 1538, 1538, 2048, 2048, 0),
		(drawing, 1539, 1539, 2048, 2048, 0),
		(drawing, 1540, 1540, 2048, 2048, 0),
		(drawing, 1541, 1541, 2048, 2048, 0),
		(drawing, 1542, 1542, 2048, 2048, 0),
		(drawing, 1543, 1543, 2048, 2048, 0),
		(drawing, 1544, 1544, 2048, 2048, 0),
		(drawing, 1545, 1545, 2048, 2048, 0),
		(drawing, 1546, 1546, 2048, 2048, 0),
		(drawing, 1547, 1547, 2048, 2048, 0),
		(drawing, 1548, 1548, 2048, 2048, 0),
		(drawing, 1549, 1549, 2048, 2048, 0),
		(drawing, 1550, 1550, 2048, 2048, 0),
		(drawing, 1551, 1551, 2048, 2048, 0),
		(drawing, 1552, 1552, 2048, 2048, 0),
		(drawing, 1553, 1553, 2048, 2048, 0),
		(drawing, 1554, 1554, 2048, 2048, 0),
		(drawing, 1555, 1555, 2048, 2048, 0),
		(drawing, 1556, 1556, 2048, 2048, 0),
		(drawing, 1557, 1557, 2048, 2048, 0),
		(drawing, 1558, 1558, 2048, 2048, 0),
		(drawing, 1559, 1559, 2048, 2048, 0),
		(drawing, 1560, 1560, 2048, 2048, 0),
		(drawing, 1561, 1561, 2048, 2048, 0),
		(drawing, 1562, 1562, 2048, 2048, 0),
		(drawing, 1563, 1563, 2048, 2048, 0),
		(drawing, 1564, 1564, 2048, 2048, 0),
		(drawing, 1565, 1565, 2048, 2048, 0),
		(drawing, 1566, 1566, 2048, 2048, 0),
		(drawing, 1567, 1567, 2048, 2048, 0),
		(drawing, 1568, 1568, 2048, 2048, 0),
		(drawing, 1569, 1569, 2048, 2048, 0),
		(drawing, 1570, 1570, 2048, 2048, 0),
		(drawing, 1571, 1571, 2048, 2048, 0),
		(drawing, 1572, 1572, 2048, 2048, 0),
		(drawing, 1573, 1573, 2048, 2048, 0),
		(drawing, 1574, 1574, 2048, 2048, 0),
		(drawing, 1575, 1575, 2048, 2048, 0),
		(drawing, 1576, 1576, 2048, 2048, 0),
		(drawing, 1577, 1577, 2048, 2048, 0),
		(drawing, 1578, 1578, 2048, 2048, 0),
		(drawing, 1579, 1579, 2048, 2048, 0),
		(drawing, 1580, 1580, 2048, 2048, 0),
		(drawing, 1581, 1581, 2048, 2048, 0),
		(drawing, 1582, 1582, 2048, 2048, 0),
		(drawing, 1583, 1583, 2048, 2048, 0),
		(drawing, 1584, 1584, 2048, 2048, 0),
		(drawing, 1585, 1585, 2048, 2048, 0),
		(drawing, 1586, 1586, 2048, 2048, 0),
		(drawing, 1587, 1587, 2048, 2048, 0),
		(drawing, 1588, 1588, 2048, 2048, 0),
		(drawing, 1589, 1589, 2048, 2048, 0),
		(drawing, 1590, 1590, 2048, 2048, 0),
		(drawing, 1591, 1591, 2048, 2048, 0),
		(drawing, 1592, 1592, 2048, 2048, 0),
		(drawing, 1593, 1593, 2048, 2048, 0),
		(drawing, 1594, 1594, 2048, 2048, 0),
		(drawing, 1595, 1595, 2048, 2048, 0),
		(drawing, 1596, 1596, 2048, 2048, 0),
		(drawing, 1597, 1597, 2048, 2048, 0),
		(drawing, 1598, 1598, 2048, 2048, 0),
		(drawing, 1599, 1599, 2048, 2048, 0),
		(drawing, 1600, 1600, 2048, 2048, 0),
		(drawing, 1601, 1601, 2048, 2048, 0),
		(drawing, 1602, 1602, 2048, 2048, 0),
		(drawing, 1603, 1603, 2048, 2048, 0),
		(drawing, 1604, 1604, 2048, 2048, 0),
		(drawing, 1605, 1605, 2048, 2048, 0),
		(drawing, 1606, 1606, 2048, 2048, 0),
		(drawing, 1607, 1607, 2048, 2048, 0),
		(drawing, 1608, 1608, 2048, 2048, 0),
		(drawing, 1609, 1609, 2048, 2048, 0),
		(drawing, 1610, 1610, 2048, 2048, 0),
		(drawing, 1611, 1611, 2048, 2048, 0),
		(drawing, 1612, 1612, 2048, 2048, 0),
		(drawing, 1613, 1613, 2048, 2048, 0),
		(drawing, 1614, 1614, 2048, 2048, 0),
		(drawing, 1615, 1615, 2048, 2048, 0),
		(drawing, 1616, 1616, 2048, 2048, 0),
		(drawing, 1617, 1617, 2048, 2048, 0),
		(drawing, 1618, 1618, 2048, 2048, 0),
		(drawing, 1619, 1619, 2048, 2048, 0),
		(drawing, 1620, 1620, 2048, 2048, 0),
		(drawing, 1621, 1621, 2048, 2048, 0),
		(drawing, 1622, 1622, 2048, 2048, 0),
		(drawing, 1623, 1623, 2048, 2048, 0),
		(drawing, 1624, 1624, 2048, 2048, 0),
		(drawing, 1625, 1625, 2048, 2048, 0),
		(drawing, 1626, 1626, 2048, 2048, 0),
		(drawing, 1627, 1627, 2048, 2048, 0),
		(drawing, 1628, 1628, 2048, 2048, 0),
		(drawing, 1629, 1629, 2048, 2048, 0),
		(drawing, 1630, 1630, 2048, 2048, 0),
		(drawing, 1631, 1631, 2048, 2048, 0),
		(drawing, 1632, 1632, 2048, 2048, 0),
		(drawing, 1633, 1633, 2048, 2048, 0),
		(drawing, 1634, 1634, 2048, 2048, 0),
		(drawing, 1635, 1635, 2048, 2048, 0),
		(drawing, 1636, 1636, 2048, 2048, 0),
		(drawing, 1637, 1637, 2048, 2048, 0),
		(drawing, 1638, 1638, 2048, 2048, 0),
		(drawing, 1639, 1639, 2048, 2048, 0),
		(drawing, 1640, 1640, 2048, 2048, 0),
		(drawing, 1641, 1641, 2048, 2048, 0),
		(drawing, 1642, 1642, 2048, 2048, 0),
		(drawing, 1643, 1643, 2048, 2048, 0),
		(drawing, 1644, 1644, 2048, 2048, 0),
		(drawing, 1645, 1645, 2048, 2048, 0),
		(drawing, 1646, 1646, 2048, 2048, 0),
		(drawing, 1647, 1647, 2048, 2048, 0),
		(drawing, 1648, 1648, 2048, 2048, 0),
		(drawing, 1649, 1649, 2048, 2048, 0),
		(drawing, 1650, 1650, 2048, 2048, 0),
		(drawing, 1651, 1651, 2048, 2048, 0),
		(drawing, 1652, 1652, 2048, 2048, 0),
		(drawing, 1653, 1653, 2048, 2048, 0),
		(drawing, 1654, 1654, 2048, 2048, 0),
		(drawing, 1655, 1655, 2048, 2048, 0),
		(drawing, 1656, 1656, 2048, 2048, 0),
		(drawing, 1657, 1657, 2048, 2048, 0),
		(drawing, 1658, 1658, 2048, 2048, 0),
		(drawing, 1659, 1659, 2048, 2048, 0),
		(drawing, 1660, 1660, 2048, 2048, 0),
		(drawing, 1661, 1661, 2048, 2048, 0),
		(drawing, 1662, 1662, 2048, 2048, 0),
		(drawing, 1663, 1663, 2048, 2048, 0),
		(drawing, 1664, 1664, 2048, 2048, 0),
		(drawing, 1665, 1665, 2048, 2048, 0),
		(drawing, 1666, 1666, 2048, 2048, 0),
		(drawing, 1667, 1667, 2048, 2048, 0),
		(drawing, 1668, 1668, 2048, 2048, 0),
		(drawing, 1669, 1669, 2048, 2048, 0),
		(drawing, 1670, 1670, 2048, 2048, 0),
		(drawing, 1671, 1671, 2048, 2048, 0),
		(drawing, 1672, 1672, 2048, 2048, 0),
		(drawing, 1673, 1673, 2048, 2048, 0),
		(drawing, 1674, 1674, 2048, 2048, 0),
		(drawing, 1675, 1675, 2048, 2048, 0),
		(drawing, 1676, 1676, 2048, 2048, 0),
		(drawing, 1677, 1677, 2048, 2048, 0),
		(drawing, 1678, 1678, 2048, 2048, 0),
		(drawing, 1679, 1679, 2048, 2048, 0),
		(drawing, 1680, 1680, 2048, 2048, 0),
		(drawing, 1681, 1681, 2048, 2048, 0),
		(drawing, 1682, 1682, 2048, 2048, 0),
		(drawing, 1683, 1683, 2048, 2048, 0),
		(drawing, 1684, 1684, 2048, 2048, 0),
		(drawing, 1685, 1685, 2048, 2048, 0),
		(drawing, 1686, 1686, 2048, 2048, 0),
		(drawing, 1687, 1687, 2048, 2048, 0),
		(drawing, 1688, 1688, 2048, 2048, 0),
		(drawing, 1689, 1689, 2048, 2048, 0),
		(drawing, 1690, 1690, 2048, 2048, 0),
		(drawing, 1691, 1691, 2048, 2048, 0),
		(drawing, 1692, 1692, 2048, 2048, 0),
		(drawing, 1693, 1693, 2048, 2048, 0),
		(drawing, 1694, 1694, 2048, 2048, 0),
		(drawing, 1695, 1695, 2048, 2048, 0),
		(drawing, 1696, 1696, 2048, 2048, 0),
		(drawing, 1697, 1697, 2048, 2048, 0),
		(drawing, 1698, 1698, 2048, 2048, 0),
		(drawing, 1699, 1699, 2048, 2048, 0),
		(drawing, 1700, 1700, 2048, 2048, 0),
		(drawing, 1701, 1701, 2048, 2048, 0),
		(drawing, 1702, 1702, 2048, 2048, 0),
		(drawing, 1703, 1703, 2048, 2048, 0),
		(drawing, 1704, 1704, 2048, 2048, 0),
		(drawing, 1705, 1705, 2048, 2048, 0),
		(drawing, 1706, 1706, 2048, 2048, 0),
		(drawing, 1707, 1707, 2048, 2048, 0),
		(drawing, 1708, 1708, 2048, 2048, 0),
		(drawing, 1709, 1709, 2048, 2048, 0),
		(drawing, 1710, 1710, 2048, 2048, 0),
		(drawing, 1711, 1711, 2048, 2048, 0),
		(drawing, 1712, 1712, 2048, 2048, 0),
		(drawing, 1713, 1713, 2048, 2048, 0),
		(drawing, 1714, 1714, 2048, 2048, 0),
		(drawing, 1715, 1715, 2048, 2048, 0),
		(drawing, 1716, 1716, 2048, 2048, 0),
		(drawing, 1717, 1717, 2048, 2048, 0),
		(drawing, 1718, 1718, 2048, 2048, 0),
		(drawing, 1719, 1719, 2048, 2048, 0),
		(drawing, 1720, 1720, 2048, 2048, 0),
		(drawing, 1721, 1721, 2048, 2048, 0),
		(drawing, 1722, 1722, 2048, 2048, 0),
		(drawing, 1723, 1723, 2048, 2048, 0),
		(drawing, 1724, 1724, 2048, 2048, 0),
		(drawing, 1725, 1725, 2048, 2048, 0),
		(drawing, 1726, 1726, 2048, 2048, 0),
		(drawing, 1727, 1727, 2048, 2048, 0),
		(drawing, 1728, 1728, 2048, 2048, 0),
		(drawing, 1729, 1729, 2048, 2048, 0),
		(drawing, 1730, 1730, 2048, 2048, 0),
		(drawing, 1731, 1731, 2048, 2048, 0),
		(drawing, 1732, 1732, 2048, 2048, 0),
		(drawing, 1733, 1733, 2048, 2048, 0),
		(drawing, 1734, 1734, 2048, 2048, 0),
		(drawing, 1735, 1735, 2048, 2048, 0),
		(drawing, 1736, 1736, 2048, 2048, 0),
		(drawing, 1737, 1737, 2048, 2048, 0),
		(drawing, 1738, 1738, 2048, 2048, 0),
		(drawing, 1739, 1739, 2048, 2048, 0),
		(drawing, 1740, 1740, 2048, 2048, 0),
		(drawing, 1741, 1741, 2048, 2048, 0),
		(drawing, 1742, 1742, 2048, 2048, 0),
		(drawing, 1743, 1743, 2048, 2048, 0),
		(drawing, 1744, 1744, 2048, 2048, 0),
		(drawing, 1745, 1745, 2048, 2048, 0),
		(drawing, 1746, 1746, 2048, 2048, 0),
		(drawing, 1747, 1747, 2048, 2048, 0),
		(drawing, 1748, 1748, 2048, 2048, 0),
		(drawing, 1749, 1749, 2048, 2048, 0),
		(drawing, 1750, 1750, 2048, 2048, 0),
		(drawing, 1751, 1751, 2048, 2048, 0),
		(drawing, 1752, 1752, 2048, 2048, 0),
		(drawing, 1753, 1753, 2048, 2048, 0),
		(drawing, 1754, 1754, 2048, 2048, 0),
		(drawing, 1755, 1755, 2048, 2048, 0),
		(drawing, 1756, 1756, 2048, 2048, 0),
		(drawing, 1757, 1757, 2048, 2048, 0),
		(drawing, 1758, 1758, 2048, 2048, 0),
		(drawing, 1759, 1759, 2048, 2048, 0),
		(drawing, 1760, 1760, 2048, 2048, 0),
		(drawing, 1761, 1761, 2048, 2048, 0),
		(drawing, 1762, 1762, 2048, 2048, 0),
		(drawing, 1763, 1763, 2048, 2048, 0),
		(drawing, 1764, 1764, 2048, 2048, 0),
		(drawing, 1765, 1765, 2048, 2048, 0),
		(drawing, 1766, 1766, 2048, 2048, 0),
		(drawing, 1767, 1767, 2048, 2048, 0),
		(drawing, 1768, 1768, 2048, 2048, 0),
		(drawing, 1769, 1769, 2048, 2048, 0),
		(drawing, 1770, 1770, 2048, 2048, 0),
		(drawing, 1771, 1771, 2048, 2048, 0),
		(drawing, 1772, 1772, 2048, 2048, 0),
		(drawing, 1773, 1773, 2048, 2048, 0),
		(drawing, 1774, 1774, 2048, 2048, 0),
		(drawing, 1775, 1775, 2048, 2048, 0),
		(drawing, 1776, 1776, 2048, 2048, 0),
		(drawing, 1777, 1777, 2048, 2048, 0),
		(drawing, 1778, 1778, 2048, 2048, 0),
		(drawing, 1779, 1779, 2048, 2048, 0),
		(drawing, 1780, 1780, 2048, 2048, 0),
		(drawing, 1781, 1781, 2048, 2048, 0),
		(drawing, 1782, 1782, 2048, 2048, 0),
		(drawing, 1783, 1783, 2048, 2048, 0),
		(drawing, 1784, 1784, 2048, 2048, 0),
		(drawing, 1785, 1785, 2048, 2048, 0),
		(drawing, 1786, 1786, 2048, 2048, 0),
		(drawing, 1787, 1787, 2048, 2048, 0),
		(drawing, 1788, 1788, 2048, 2048, 0),
		(drawing, 1789, 1789, 2048, 2048, 0),
		(drawing, 1790, 1790, 2048, 2048, 0),
		(drawing, 1791, 1791, 2048, 2048, 0),
		(drawing, 1792, 1792, 2048, 2048, 0),
		(drawing, 1793, 1793, 2048, 2048, 0),
		(drawing, 1794, 1794, 2048, 2048, 0),
		(drawing, 1795, 1795, 2048, 2048, 0),
		(drawing, 1796, 1796, 2048, 2048, 0),
		(drawing, 1797, 1797, 2048, 2048, 0),
		(drawing, 1798, 1798, 2048, 2048, 0),
		(drawing, 1799, 1799, 2048, 2048, 0),
		(drawing, 1800, 1800, 2048, 2048, 0),
		(drawing, 1801, 1801, 2048, 2048, 0),
		(drawing, 1802, 1802, 2048, 2048, 0),
		(drawing, 1803, 1803, 2048, 2048, 0),
		(drawing, 1804, 1804, 2048, 2048, 0),
		(drawing, 1805, 1805, 2048, 2048, 0),
		(drawing, 1806, 1806, 2048, 2048, 0),
		(drawing, 1807, 1807, 2048, 2048, 0),
		(drawing, 1808, 1808, 2048, 2048, 0),
		(drawing, 1809, 1809, 2048, 2048, 0),
		(drawing, 1810, 1810, 2048, 2048, 0),
		(drawing, 1811, 1811, 2048, 2048, 0),
		(drawing, 1812, 1812, 2048, 2048, 0),
		(drawing, 1813, 1813, 2048, 2048, 0),
		(drawing, 1814, 1814, 2048, 2048, 0),
		(drawing, 1815, 1815, 2048, 2048, 0),
		(drawing, 1816, 1816, 2048, 2048, 0),
		(drawing, 1817, 1817, 2048, 2048, 0),
		(drawing, 1818, 1818, 2048, 2048, 0),
		(drawing, 1819, 1819, 2048, 2048, 0),
		(drawing, 1820, 1820, 2048, 2048, 0),
		(drawing, 1821, 1821, 2048, 2048, 0),
		(drawing, 1822, 1822, 2048, 2048, 0),
		(drawing, 1823, 1823, 2048, 2048, 0),
		(drawing, 1824, 1824, 2048, 2048, 0),
		(drawing, 1825, 1825, 2048, 2048, 0),
		(drawing, 1826, 1826, 2048, 2048, 0),
		(drawing, 1827, 1827, 2048, 2048, 0),
		(drawing, 1828, 1828, 2048, 2048, 0),
		(drawing, 1829, 1829, 2048, 2048, 0),
		(drawing, 1830, 1830, 2048, 2048, 0),
		(drawing, 1831, 1831, 2048, 2048, 0),
		(drawing, 1832, 1832, 2048, 2048, 0),
		(drawing, 1833, 1833, 2048, 2048, 0),
		(drawing, 1834, 1834, 2048, 2048, 0),
		(drawing, 1835, 1835, 2048, 2048, 0),
		(drawing, 1836, 1836, 2048, 2048, 0),
		(drawing, 1837, 1837, 2048, 2048, 0),
		(drawing, 1838, 1838, 2048, 2048, 0),
		(drawing, 1839, 1839, 2048, 2048, 0),
		(drawing, 1840, 1840, 2048, 2048, 0),
		(drawing, 1841, 1841, 2048, 2048, 0),
		(drawing, 1842, 1842, 2048, 2048, 0),
		(drawing, 1843, 1843, 2048, 2048, 0),
		(drawing, 1844, 1844, 2048, 2048, 0),
		(drawing, 1845, 1845, 2048, 2048, 0),
		(drawing, 1846, 1846, 2048, 2048, 0),
		(drawing, 1847, 1847, 2048, 2048, 0),
		(drawing, 1848, 1848, 2048, 2048, 0),
		(drawing, 1849, 1849, 2048, 2048, 0),
		(drawing, 1850, 1850, 2048, 2048, 0),
		(drawing, 1851, 1851, 2048, 2048, 0),
		(drawing, 1852, 1852, 2048, 2048, 0),
		(drawing, 1853, 1853, 2048, 2048, 0),
		(drawing, 1854, 1854, 2048, 2048, 0),
		(drawing, 1855, 1855, 2048, 2048, 0),
		(drawing, 1856, 1856, 2048, 2048, 0),
		(drawing, 1857, 1857, 2048, 2048, 0),
		(drawing, 1858, 1858, 2048, 2048, 0),
		(drawing, 1859, 1859, 2048, 2048, 0),
		(drawing, 1860, 1860, 2048, 2048, 0),
		(drawing, 1861, 1861, 2048, 2048, 0),
		(drawing, 1862, 1862, 2048, 2048, 0),
		(drawing, 1863, 1863, 2048, 2048, 0),
		(drawing, 1864, 1864, 2048, 2048, 0),
		(drawing, 1865, 1865, 2048, 2048, 0),
		(drawing, 1866, 1866, 2048, 2048, 0),
		(drawing, 1867, 1867, 2048, 2048, 0),
		(drawing, 1868, 1868, 2048, 2048, 0),
		(drawing, 1869, 1869, 2048, 2048, 0),
		(drawing, 1870, 1870, 2048, 2048, 0),
		(drawing, 1871, 1871, 2048, 2048, 0),
		(drawing, 1872, 1872, 2048, 2048, 0),
		(drawing, 1873, 1873, 2048, 2048, 0),
		(drawing, 1874, 1874, 2048, 2048, 0),
		(drawing, 1875, 1875, 2048, 2048, 0),
		(drawing, 1876, 1876, 2048, 2048, 0),
		(drawing, 1877, 1877, 2048, 2048, 0),
		(drawing, 1878, 1878, 2048, 2048, 0),
		(drawing, 1879, 1879, 2048, 2048, 0),
		(drawing, 1880, 1880, 2048, 2048, 0),
		(drawing, 1881, 1881, 2048, 2048, 0),
		(drawing, 1882, 1882, 2048, 2048, 0),
		(drawing, 1883, 1883, 2048, 2048, 0),
		(drawing, 1884, 1884, 2048, 2048, 0),
		(drawing, 1885, 1885, 2048, 2048, 0),
		(drawing, 1886, 1886, 2048, 2048, 0),
		(drawing, 1887, 1887, 2048, 2048, 0),
		(drawing, 1888, 1888, 2048, 2048, 0),
		(drawing, 1889, 1889, 2048, 2048, 0),
		(drawing, 1890, 1890, 2048, 2048, 0),
		(drawing, 1891, 1891, 2048, 2048, 0),
		(drawing, 1892, 1892, 2048, 2048, 0),
		(drawing, 1893, 1893, 2048, 2048, 0),
		(drawing, 1894, 1894, 2048, 2048, 0),
		(drawing, 1895, 1895, 2048, 2048, 0),
		(drawing, 1896, 1896, 2048, 2048, 0),
		(drawing, 1897, 1897, 2048, 2048, 0),
		(drawing, 1898, 1898, 2048, 2048, 0),
		(drawing, 1899, 1899, 2048, 2048, 0),
		(drawing, 1900, 1900, 2048, 2048, 0),
		(drawing, 1901, 1901, 2048, 2048, 0),
		(drawing, 1902, 1902, 2048, 2048, 0),
		(drawing, 1903, 1903, 2048, 2048, 0),
		(drawing, 1904, 1904, 2048, 2048, 0),
		(drawing, 1905, 1905, 2048, 2048, 0),
		(drawing, 1906, 1906, 2048, 2048, 0),
		(drawing, 1907, 1907, 2048, 2048, 0),
		(drawing, 1908, 1908, 2048, 2048, 0),
		(drawing, 1909, 1909, 2048, 2048, 0),
		(drawing, 1910, 1910, 2048, 2048, 0),
		(drawing, 1911, 1911, 2048, 2048, 0),
		(drawing, 1912, 1912, 2048, 2048, 0),
		(drawing, 1913, 1913, 2048, 2048, 0),
		(drawing, 1914, 1914, 2048, 2048, 0),
		(drawing, 1915, 1915, 2048, 2048, 0),
		(drawing, 1916, 1916, 2048, 2048, 0),
		(drawing, 1917, 1917, 2048, 2048, 0),
		(drawing, 1918, 1918, 2048, 2048, 0),
		(drawing, 1919, 1919, 2048, 2048, 0),
		(drawing, 1920, 1920, 2048, 2048, 0),
		(drawing, 1921, 1921, 2048, 2048, 0),
		(drawing, 1922, 1922, 2048, 2048, 0),
		(drawing, 1923, 1923, 2048, 2048, 0),
		(drawing, 1924, 1924, 2048, 2048, 0),
		(drawing, 1925, 1925, 2048, 2048, 0),
		(drawing, 1926, 1926, 2048, 2048, 0),
		(drawing, 1927, 1927, 2048, 2048, 0),
		(drawing, 1928, 1928, 2048, 2048, 0),
		(drawing, 1929, 1929, 2048, 2048, 0),
		(drawing, 1930, 1930, 2048, 2048, 0),
		(drawing, 1931, 1931, 2048, 2048, 0),
		(drawing, 1932, 1932, 2048, 2048, 0),
		(drawing, 1933, 1933, 2048, 2048, 0),
		(drawing, 1934, 1934, 2048, 2048, 0),
		(drawing, 1935, 1935, 2048, 2048, 0),
		(drawing, 1936, 1936, 2048, 2048, 0),
		(drawing, 1937, 1937, 2048, 2048, 0),
		(drawing, 1938, 1938, 2048, 2048, 0),
		(drawing, 1939, 1939, 2048, 2048, 0),
		(drawing, 1940, 1940, 2048, 2048, 0),
		(drawing, 1941, 1941, 2048, 2048, 0),
		(drawing, 1942, 1942, 2048, 2048, 0),
		(drawing, 1943, 1943, 2048, 2048, 0),
		(drawing, 1944, 1944, 2048, 2048, 0),
		(drawing, 1945, 1945, 2048, 2048, 0),
		(drawing, 1946, 1946, 2048, 2048, 0),
		(drawing, 1947, 1947, 2048, 2048, 0),
		(drawing, 1948, 1948, 2048, 2048, 0),
		(drawing, 1949, 1949, 2048, 2048, 0),
		(drawing, 1950, 1950, 2048, 2048, 0),
		(drawing, 1951, 1951, 2048, 2048, 0),
		(drawing, 1952, 1952, 2048, 2048, 0),
		(drawing, 1953, 1953, 2048, 2048, 0),
		(drawing, 1954, 1954, 2048, 2048, 0),
		(drawing, 1955, 1955, 2048, 2048, 0),
		(drawing, 1956, 1956, 2048, 2048, 0),
		(drawing, 1957, 1957, 2048, 2048, 0),
		(drawing, 1958, 1958, 2048, 2048, 0),
		(drawing, 1959, 1959, 2048, 2048, 0),
		(drawing, 1960, 1960, 2048, 2048, 0),
		(drawing, 1961, 1961, 2048, 2048, 0),
		(drawing, 1962, 1962, 2048, 2048, 0),
		(drawing, 1963, 1963, 2048, 2048, 0),
		(drawing, 1964, 1964, 2048, 2048, 0),
		(drawing, 1965, 1965, 2048, 2048, 0),
		(drawing, 1966, 1966, 2048, 2048, 0),
		(drawing, 1967, 1967, 2048, 2048, 0),
		(drawing, 1968, 1968, 2048, 2048, 0),
		(drawing, 1969, 1969, 2048, 2048, 0),
		(drawing, 1970, 1970, 2048, 2048, 0),
		(drawing, 1971, 1971, 2048, 2048, 0),
		(drawing, 1972, 1972, 2048, 2048, 0),
		(drawing, 1973, 1973, 2048, 2048, 0),
		(drawing, 1974, 1974, 2048, 2048, 0),
		(drawing, 1975, 1975, 2048, 2048, 0),
		(drawing, 1976, 1976, 2048, 2048, 0),
		(drawing, 1977, 1977, 2048, 2048, 0),
		(drawing, 1978, 1978, 2048, 2048, 0),
		(drawing, 1979, 1979, 2048, 2048, 0),
		(drawing, 1980, 1980, 2048, 2048, 0),
		(drawing, 1981, 1981, 2048, 2048, 0),
		(drawing, 1982, 1982, 2048, 2048, 0),
		(drawing, 1983, 1983, 2048, 2048, 0),
		(drawing, 1984, 1984, 2048, 2048, 0),
		(drawing, 1985, 1985, 2048, 2048, 0),
		(drawing, 1986, 1986, 2048, 2048, 0),
		(drawing, 1987, 1987, 2048, 2048, 0),
		(drawing, 1988, 1988, 2048, 2048, 0),
		(drawing, 1989, 1989, 2048, 2048, 0),
		(drawing, 1990, 1990, 2048, 2048, 0),
		(drawing, 1991, 1991, 2048, 2048, 0),
		(drawing, 1992, 1992, 2048, 2048, 0),
		(drawing, 1993, 1993, 2048, 2048, 0),
		(drawing, 1994, 1994, 2048, 2048, 0),
		(drawing, 1995, 1995, 2048, 2048, 0),
		(drawing, 1996, 1996, 2048, 2048, 0),
		(drawing, 1997, 1997, 2048, 2048, 0),
		(drawing, 1998, 1998, 2048, 2048, 0),
		(drawing, 1999, 1999, 2048, 2048, 0),
		(drawing, 2000, 2000, 2048, 2048, 0),
		(drawing, 2001, 2001, 2048, 2048, 0),
		(drawing, 2002, 2002, 2048, 2048, 0),
		(drawing, 2003, 2003, 2048, 2048, 0),
		(drawing, 2004, 2004, 2048, 2048, 0),
		(drawing, 2005, 2005, 2048, 2048, 0),
		(drawing, 2006, 2006, 2048, 2048, 0),
		(drawing, 2007, 2007, 2048, 2048, 0),
		(drawing, 2008, 2008, 2048, 2048, 0),
		(drawing, 2009, 2009, 2048, 2048, 0),
		(drawing, 2010, 2010, 2048, 2048, 0),
		(drawing, 2011, 2011, 2048, 2048, 0),
		(drawing, 2012, 2012, 2048, 2048, 0),
		(drawing, 2013, 2013, 2048, 2048, 0),
		(drawing, 2014, 2014, 2048, 2048, 0),
		(drawing, 2015, 2015, 2048, 2048, 0),
		(drawing, 2016, 2016, 2048, 2048, 0),
		(drawing, 2017, 2017, 2048, 2048, 0),
		(drawing, 2018, 2018, 2048, 2048, 0),
		(drawing, 2019, 2019, 2048, 2048, 0),
		(drawing, 2020, 2020, 2048, 2048, 0),
		(drawing, 2021, 2021, 2048, 2048, 0),
		(drawing, 2022, 2022, 2048, 2048, 0),
		(drawing, 2023, 2023, 2048, 2048, 0),
		(drawing, 2024, 2024, 2048, 2048, 0),
		(drawing, 2025, 2025, 2048, 2048, 0),
		(drawing, 2026, 2026, 2048, 2048, 0),
		(drawing, 2027, 2027, 2048, 2048, 0),
		(drawing, 2028, 2028, 2048, 2048, 0),
		(drawing, 2029, 2029, 2048, 2048, 0),
		(drawing, 2030, 2030, 2048, 2048, 0),
		(drawing, 2031, 2031, 2048, 2048, 0),
		(drawing, 2032, 2032, 2048, 2048, 0),
		(drawing, 2033, 2033, 2048, 2048, 0),
		(drawing, 2034, 2034, 2048, 2048, 0),
		(drawing, 2035, 2035, 2048, 2048, 0),
		(drawing, 2036, 2036, 2048, 2048, 0),
		(drawing, 2037, 2037, 2048, 2048, 0),
		(drawing, 2038, 2038, 2048, 2048, 0),
		(drawing, 2039, 2039, 2048, 2048, 0),
		(drawing, 2040, 2040, 2048, 2048, 0),
		(drawing, 2041, 2041, 2048, 2048, 0),
		(drawing, 2042, 2042, 2048, 2048, 0),
		(drawing, 2043, 2043, 2048, 2048, 0),
		(drawing, 2044, 2044, 2048, 2048, 0),
		(drawing, 2045, 2045, 2048, 2048, 0),
		(drawing, 2046, 2046, 2048, 2048, 0),
		(drawing, 2047, 2047, 2048, 2048, 0),
		(done, 2048, 2048, 2048, 2048, 0)
	);
END PACKAGE ex1_data_pak;
