-- advanced test 4
-- draw line from (0,0) to (4095,4095)
-- NOTE * xin,yin are 12bits logic vectors
--------* the maximum value of them is b1111,1111,1111 which is 4095 in decimal
--------* this test is for the case of maximum possible value of xin,yin

PACKAGE ex1_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 0, 0, 0),
		(start, 0, 0, 4095, 4095, 0),
		(drawing, 0, 0, 4095, 4095, 0),
		(drawing, 1, 1, 4095, 4095, 0),
		(drawing, 2, 2, 4095, 4095, 0),
		(drawing, 3, 3, 4095, 4095, 0),
		(drawing, 4, 4, 4095, 4095, 0),
		(drawing, 5, 5, 4095, 4095, 0),
		(drawing, 6, 6, 4095, 4095, 0),
		(drawing, 7, 7, 4095, 4095, 0),
		(drawing, 8, 8, 4095, 4095, 0),
		(drawing, 9, 9, 4095, 4095, 0),
		(drawing, 10, 10, 4095, 4095, 0),
		(drawing, 11, 11, 4095, 4095, 0),
		(drawing, 12, 12, 4095, 4095, 0),
		(drawing, 13, 13, 4095, 4095, 0),
		(drawing, 14, 14, 4095, 4095, 0),
		(drawing, 15, 15, 4095, 4095, 0),
		(drawing, 16, 16, 4095, 4095, 0),
		(drawing, 17, 17, 4095, 4095, 0),
		(drawing, 18, 18, 4095, 4095, 0),
		(drawing, 19, 19, 4095, 4095, 0),
		(drawing, 20, 20, 4095, 4095, 0),
		(drawing, 21, 21, 4095, 4095, 0),
		(drawing, 22, 22, 4095, 4095, 0),
		(drawing, 23, 23, 4095, 4095, 0),
		(drawing, 24, 24, 4095, 4095, 0),
		(drawing, 25, 25, 4095, 4095, 0),
		(drawing, 26, 26, 4095, 4095, 0),
		(drawing, 27, 27, 4095, 4095, 0),
		(drawing, 28, 28, 4095, 4095, 0),
		(drawing, 29, 29, 4095, 4095, 0),
		(drawing, 30, 30, 4095, 4095, 0),
		(drawing, 31, 31, 4095, 4095, 0),
		(drawing, 32, 32, 4095, 4095, 0),
		(drawing, 33, 33, 4095, 4095, 0),
		(drawing, 34, 34, 4095, 4095, 0),
		(drawing, 35, 35, 4095, 4095, 0),
		(drawing, 36, 36, 4095, 4095, 0),
		(drawing, 37, 37, 4095, 4095, 0),
		(drawing, 38, 38, 4095, 4095, 0),
		(drawing, 39, 39, 4095, 4095, 0),
		(drawing, 40, 40, 4095, 4095, 0),
		(drawing, 41, 41, 4095, 4095, 0),
		(drawing, 42, 42, 4095, 4095, 0),
		(drawing, 43, 43, 4095, 4095, 0),
		(drawing, 44, 44, 4095, 4095, 0),
		(drawing, 45, 45, 4095, 4095, 0),
		(drawing, 46, 46, 4095, 4095, 0),
		(drawing, 47, 47, 4095, 4095, 0),
		(drawing, 48, 48, 4095, 4095, 0),
		(drawing, 49, 49, 4095, 4095, 0),
		(drawing, 50, 50, 4095, 4095, 0),
		(drawing, 51, 51, 4095, 4095, 0),
		(drawing, 52, 52, 4095, 4095, 0),
		(drawing, 53, 53, 4095, 4095, 0),
		(drawing, 54, 54, 4095, 4095, 0),
		(drawing, 55, 55, 4095, 4095, 0),
		(drawing, 56, 56, 4095, 4095, 0),
		(drawing, 57, 57, 4095, 4095, 0),
		(drawing, 58, 58, 4095, 4095, 0),
		(drawing, 59, 59, 4095, 4095, 0),
		(drawing, 60, 60, 4095, 4095, 0),
		(drawing, 61, 61, 4095, 4095, 0),
		(drawing, 62, 62, 4095, 4095, 0),
		(drawing, 63, 63, 4095, 4095, 0),
		(drawing, 64, 64, 4095, 4095, 0),
		(drawing, 65, 65, 4095, 4095, 0),
		(drawing, 66, 66, 4095, 4095, 0),
		(drawing, 67, 67, 4095, 4095, 0),
		(drawing, 68, 68, 4095, 4095, 0),
		(drawing, 69, 69, 4095, 4095, 0),
		(drawing, 70, 70, 4095, 4095, 0),
		(drawing, 71, 71, 4095, 4095, 0),
		(drawing, 72, 72, 4095, 4095, 0),
		(drawing, 73, 73, 4095, 4095, 0),
		(drawing, 74, 74, 4095, 4095, 0),
		(drawing, 75, 75, 4095, 4095, 0),
		(drawing, 76, 76, 4095, 4095, 0),
		(drawing, 77, 77, 4095, 4095, 0),
		(drawing, 78, 78, 4095, 4095, 0),
		(drawing, 79, 79, 4095, 4095, 0),
		(drawing, 80, 80, 4095, 4095, 0),
		(drawing, 81, 81, 4095, 4095, 0),
		(drawing, 82, 82, 4095, 4095, 0),
		(drawing, 83, 83, 4095, 4095, 0),
		(drawing, 84, 84, 4095, 4095, 0),
		(drawing, 85, 85, 4095, 4095, 0),
		(drawing, 86, 86, 4095, 4095, 0),
		(drawing, 87, 87, 4095, 4095, 0),
		(drawing, 88, 88, 4095, 4095, 0),
		(drawing, 89, 89, 4095, 4095, 0),
		(drawing, 90, 90, 4095, 4095, 0),
		(drawing, 91, 91, 4095, 4095, 0),
		(drawing, 92, 92, 4095, 4095, 0),
		(drawing, 93, 93, 4095, 4095, 0),
		(drawing, 94, 94, 4095, 4095, 0),
		(drawing, 95, 95, 4095, 4095, 0),
		(drawing, 96, 96, 4095, 4095, 0),
		(drawing, 97, 97, 4095, 4095, 0),
		(drawing, 98, 98, 4095, 4095, 0),
		(drawing, 99, 99, 4095, 4095, 0),
		(drawing, 100, 100, 4095, 4095, 0),
		(drawing, 101, 101, 4095, 4095, 0),
		(drawing, 102, 102, 4095, 4095, 0),
		(drawing, 103, 103, 4095, 4095, 0),
		(drawing, 104, 104, 4095, 4095, 0),
		(drawing, 105, 105, 4095, 4095, 0),
		(drawing, 106, 106, 4095, 4095, 0),
		(drawing, 107, 107, 4095, 4095, 0),
		(drawing, 108, 108, 4095, 4095, 0),
		(drawing, 109, 109, 4095, 4095, 0),
		(drawing, 110, 110, 4095, 4095, 0),
		(drawing, 111, 111, 4095, 4095, 0),
		(drawing, 112, 112, 4095, 4095, 0),
		(drawing, 113, 113, 4095, 4095, 0),
		(drawing, 114, 114, 4095, 4095, 0),
		(drawing, 115, 115, 4095, 4095, 0),
		(drawing, 116, 116, 4095, 4095, 0),
		(drawing, 117, 117, 4095, 4095, 0),
		(drawing, 118, 118, 4095, 4095, 0),
		(drawing, 119, 119, 4095, 4095, 0),
		(drawing, 120, 120, 4095, 4095, 0),
		(drawing, 121, 121, 4095, 4095, 0),
		(drawing, 122, 122, 4095, 4095, 0),
		(drawing, 123, 123, 4095, 4095, 0),
		(drawing, 124, 124, 4095, 4095, 0),
		(drawing, 125, 125, 4095, 4095, 0),
		(drawing, 126, 126, 4095, 4095, 0),
		(drawing, 127, 127, 4095, 4095, 0),
		(drawing, 128, 128, 4095, 4095, 0),
		(drawing, 129, 129, 4095, 4095, 0),
		(drawing, 130, 130, 4095, 4095, 0),
		(drawing, 131, 131, 4095, 4095, 0),
		(drawing, 132, 132, 4095, 4095, 0),
		(drawing, 133, 133, 4095, 4095, 0),
		(drawing, 134, 134, 4095, 4095, 0),
		(drawing, 135, 135, 4095, 4095, 0),
		(drawing, 136, 136, 4095, 4095, 0),
		(drawing, 137, 137, 4095, 4095, 0),
		(drawing, 138, 138, 4095, 4095, 0),
		(drawing, 139, 139, 4095, 4095, 0),
		(drawing, 140, 140, 4095, 4095, 0),
		(drawing, 141, 141, 4095, 4095, 0),
		(drawing, 142, 142, 4095, 4095, 0),
		(drawing, 143, 143, 4095, 4095, 0),
		(drawing, 144, 144, 4095, 4095, 0),
		(drawing, 145, 145, 4095, 4095, 0),
		(drawing, 146, 146, 4095, 4095, 0),
		(drawing, 147, 147, 4095, 4095, 0),
		(drawing, 148, 148, 4095, 4095, 0),
		(drawing, 149, 149, 4095, 4095, 0),
		(drawing, 150, 150, 4095, 4095, 0),
		(drawing, 151, 151, 4095, 4095, 0),
		(drawing, 152, 152, 4095, 4095, 0),
		(drawing, 153, 153, 4095, 4095, 0),
		(drawing, 154, 154, 4095, 4095, 0),
		(drawing, 155, 155, 4095, 4095, 0),
		(drawing, 156, 156, 4095, 4095, 0),
		(drawing, 157, 157, 4095, 4095, 0),
		(drawing, 158, 158, 4095, 4095, 0),
		(drawing, 159, 159, 4095, 4095, 0),
		(drawing, 160, 160, 4095, 4095, 0),
		(drawing, 161, 161, 4095, 4095, 0),
		(drawing, 162, 162, 4095, 4095, 0),
		(drawing, 163, 163, 4095, 4095, 0),
		(drawing, 164, 164, 4095, 4095, 0),
		(drawing, 165, 165, 4095, 4095, 0),
		(drawing, 166, 166, 4095, 4095, 0),
		(drawing, 167, 167, 4095, 4095, 0),
		(drawing, 168, 168, 4095, 4095, 0),
		(drawing, 169, 169, 4095, 4095, 0),
		(drawing, 170, 170, 4095, 4095, 0),
		(drawing, 171, 171, 4095, 4095, 0),
		(drawing, 172, 172, 4095, 4095, 0),
		(drawing, 173, 173, 4095, 4095, 0),
		(drawing, 174, 174, 4095, 4095, 0),
		(drawing, 175, 175, 4095, 4095, 0),
		(drawing, 176, 176, 4095, 4095, 0),
		(drawing, 177, 177, 4095, 4095, 0),
		(drawing, 178, 178, 4095, 4095, 0),
		(drawing, 179, 179, 4095, 4095, 0),
		(drawing, 180, 180, 4095, 4095, 0),
		(drawing, 181, 181, 4095, 4095, 0),
		(drawing, 182, 182, 4095, 4095, 0),
		(drawing, 183, 183, 4095, 4095, 0),
		(drawing, 184, 184, 4095, 4095, 0),
		(drawing, 185, 185, 4095, 4095, 0),
		(drawing, 186, 186, 4095, 4095, 0),
		(drawing, 187, 187, 4095, 4095, 0),
		(drawing, 188, 188, 4095, 4095, 0),
		(drawing, 189, 189, 4095, 4095, 0),
		(drawing, 190, 190, 4095, 4095, 0),
		(drawing, 191, 191, 4095, 4095, 0),
		(drawing, 192, 192, 4095, 4095, 0),
		(drawing, 193, 193, 4095, 4095, 0),
		(drawing, 194, 194, 4095, 4095, 0),
		(drawing, 195, 195, 4095, 4095, 0),
		(drawing, 196, 196, 4095, 4095, 0),
		(drawing, 197, 197, 4095, 4095, 0),
		(drawing, 198, 198, 4095, 4095, 0),
		(drawing, 199, 199, 4095, 4095, 0),
		(drawing, 200, 200, 4095, 4095, 0),
		(drawing, 201, 201, 4095, 4095, 0),
		(drawing, 202, 202, 4095, 4095, 0),
		(drawing, 203, 203, 4095, 4095, 0),
		(drawing, 204, 204, 4095, 4095, 0),
		(drawing, 205, 205, 4095, 4095, 0),
		(drawing, 206, 206, 4095, 4095, 0),
		(drawing, 207, 207, 4095, 4095, 0),
		(drawing, 208, 208, 4095, 4095, 0),
		(drawing, 209, 209, 4095, 4095, 0),
		(drawing, 210, 210, 4095, 4095, 0),
		(drawing, 211, 211, 4095, 4095, 0),
		(drawing, 212, 212, 4095, 4095, 0),
		(drawing, 213, 213, 4095, 4095, 0),
		(drawing, 214, 214, 4095, 4095, 0),
		(drawing, 215, 215, 4095, 4095, 0),
		(drawing, 216, 216, 4095, 4095, 0),
		(drawing, 217, 217, 4095, 4095, 0),
		(drawing, 218, 218, 4095, 4095, 0),
		(drawing, 219, 219, 4095, 4095, 0),
		(drawing, 220, 220, 4095, 4095, 0),
		(drawing, 221, 221, 4095, 4095, 0),
		(drawing, 222, 222, 4095, 4095, 0),
		(drawing, 223, 223, 4095, 4095, 0),
		(drawing, 224, 224, 4095, 4095, 0),
		(drawing, 225, 225, 4095, 4095, 0),
		(drawing, 226, 226, 4095, 4095, 0),
		(drawing, 227, 227, 4095, 4095, 0),
		(drawing, 228, 228, 4095, 4095, 0),
		(drawing, 229, 229, 4095, 4095, 0),
		(drawing, 230, 230, 4095, 4095, 0),
		(drawing, 231, 231, 4095, 4095, 0),
		(drawing, 232, 232, 4095, 4095, 0),
		(drawing, 233, 233, 4095, 4095, 0),
		(drawing, 234, 234, 4095, 4095, 0),
		(drawing, 235, 235, 4095, 4095, 0),
		(drawing, 236, 236, 4095, 4095, 0),
		(drawing, 237, 237, 4095, 4095, 0),
		(drawing, 238, 238, 4095, 4095, 0),
		(drawing, 239, 239, 4095, 4095, 0),
		(drawing, 240, 240, 4095, 4095, 0),
		(drawing, 241, 241, 4095, 4095, 0),
		(drawing, 242, 242, 4095, 4095, 0),
		(drawing, 243, 243, 4095, 4095, 0),
		(drawing, 244, 244, 4095, 4095, 0),
		(drawing, 245, 245, 4095, 4095, 0),
		(drawing, 246, 246, 4095, 4095, 0),
		(drawing, 247, 247, 4095, 4095, 0),
		(drawing, 248, 248, 4095, 4095, 0),
		(drawing, 249, 249, 4095, 4095, 0),
		(drawing, 250, 250, 4095, 4095, 0),
		(drawing, 251, 251, 4095, 4095, 0),
		(drawing, 252, 252, 4095, 4095, 0),
		(drawing, 253, 253, 4095, 4095, 0),
		(drawing, 254, 254, 4095, 4095, 0),
		(drawing, 255, 255, 4095, 4095, 0),
		(drawing, 256, 256, 4095, 4095, 0),
		(drawing, 257, 257, 4095, 4095, 0),
		(drawing, 258, 258, 4095, 4095, 0),
		(drawing, 259, 259, 4095, 4095, 0),
		(drawing, 260, 260, 4095, 4095, 0),
		(drawing, 261, 261, 4095, 4095, 0),
		(drawing, 262, 262, 4095, 4095, 0),
		(drawing, 263, 263, 4095, 4095, 0),
		(drawing, 264, 264, 4095, 4095, 0),
		(drawing, 265, 265, 4095, 4095, 0),
		(drawing, 266, 266, 4095, 4095, 0),
		(drawing, 267, 267, 4095, 4095, 0),
		(drawing, 268, 268, 4095, 4095, 0),
		(drawing, 269, 269, 4095, 4095, 0),
		(drawing, 270, 270, 4095, 4095, 0),
		(drawing, 271, 271, 4095, 4095, 0),
		(drawing, 272, 272, 4095, 4095, 0),
		(drawing, 273, 273, 4095, 4095, 0),
		(drawing, 274, 274, 4095, 4095, 0),
		(drawing, 275, 275, 4095, 4095, 0),
		(drawing, 276, 276, 4095, 4095, 0),
		(drawing, 277, 277, 4095, 4095, 0),
		(drawing, 278, 278, 4095, 4095, 0),
		(drawing, 279, 279, 4095, 4095, 0),
		(drawing, 280, 280, 4095, 4095, 0),
		(drawing, 281, 281, 4095, 4095, 0),
		(drawing, 282, 282, 4095, 4095, 0),
		(drawing, 283, 283, 4095, 4095, 0),
		(drawing, 284, 284, 4095, 4095, 0),
		(drawing, 285, 285, 4095, 4095, 0),
		(drawing, 286, 286, 4095, 4095, 0),
		(drawing, 287, 287, 4095, 4095, 0),
		(drawing, 288, 288, 4095, 4095, 0),
		(drawing, 289, 289, 4095, 4095, 0),
		(drawing, 290, 290, 4095, 4095, 0),
		(drawing, 291, 291, 4095, 4095, 0),
		(drawing, 292, 292, 4095, 4095, 0),
		(drawing, 293, 293, 4095, 4095, 0),
		(drawing, 294, 294, 4095, 4095, 0),
		(drawing, 295, 295, 4095, 4095, 0),
		(drawing, 296, 296, 4095, 4095, 0),
		(drawing, 297, 297, 4095, 4095, 0),
		(drawing, 298, 298, 4095, 4095, 0),
		(drawing, 299, 299, 4095, 4095, 0),
		(drawing, 300, 300, 4095, 4095, 0),
		(drawing, 301, 301, 4095, 4095, 0),
		(drawing, 302, 302, 4095, 4095, 0),
		(drawing, 303, 303, 4095, 4095, 0),
		(drawing, 304, 304, 4095, 4095, 0),
		(drawing, 305, 305, 4095, 4095, 0),
		(drawing, 306, 306, 4095, 4095, 0),
		(drawing, 307, 307, 4095, 4095, 0),
		(drawing, 308, 308, 4095, 4095, 0),
		(drawing, 309, 309, 4095, 4095, 0),
		(drawing, 310, 310, 4095, 4095, 0),
		(drawing, 311, 311, 4095, 4095, 0),
		(drawing, 312, 312, 4095, 4095, 0),
		(drawing, 313, 313, 4095, 4095, 0),
		(drawing, 314, 314, 4095, 4095, 0),
		(drawing, 315, 315, 4095, 4095, 0),
		(drawing, 316, 316, 4095, 4095, 0),
		(drawing, 317, 317, 4095, 4095, 0),
		(drawing, 318, 318, 4095, 4095, 0),
		(drawing, 319, 319, 4095, 4095, 0),
		(drawing, 320, 320, 4095, 4095, 0),
		(drawing, 321, 321, 4095, 4095, 0),
		(drawing, 322, 322, 4095, 4095, 0),
		(drawing, 323, 323, 4095, 4095, 0),
		(drawing, 324, 324, 4095, 4095, 0),
		(drawing, 325, 325, 4095, 4095, 0),
		(drawing, 326, 326, 4095, 4095, 0),
		(drawing, 327, 327, 4095, 4095, 0),
		(drawing, 328, 328, 4095, 4095, 0),
		(drawing, 329, 329, 4095, 4095, 0),
		(drawing, 330, 330, 4095, 4095, 0),
		(drawing, 331, 331, 4095, 4095, 0),
		(drawing, 332, 332, 4095, 4095, 0),
		(drawing, 333, 333, 4095, 4095, 0),
		(drawing, 334, 334, 4095, 4095, 0),
		(drawing, 335, 335, 4095, 4095, 0),
		(drawing, 336, 336, 4095, 4095, 0),
		(drawing, 337, 337, 4095, 4095, 0),
		(drawing, 338, 338, 4095, 4095, 0),
		(drawing, 339, 339, 4095, 4095, 0),
		(drawing, 340, 340, 4095, 4095, 0),
		(drawing, 341, 341, 4095, 4095, 0),
		(drawing, 342, 342, 4095, 4095, 0),
		(drawing, 343, 343, 4095, 4095, 0),
		(drawing, 344, 344, 4095, 4095, 0),
		(drawing, 345, 345, 4095, 4095, 0),
		(drawing, 346, 346, 4095, 4095, 0),
		(drawing, 347, 347, 4095, 4095, 0),
		(drawing, 348, 348, 4095, 4095, 0),
		(drawing, 349, 349, 4095, 4095, 0),
		(drawing, 350, 350, 4095, 4095, 0),
		(drawing, 351, 351, 4095, 4095, 0),
		(drawing, 352, 352, 4095, 4095, 0),
		(drawing, 353, 353, 4095, 4095, 0),
		(drawing, 354, 354, 4095, 4095, 0),
		(drawing, 355, 355, 4095, 4095, 0),
		(drawing, 356, 356, 4095, 4095, 0),
		(drawing, 357, 357, 4095, 4095, 0),
		(drawing, 358, 358, 4095, 4095, 0),
		(drawing, 359, 359, 4095, 4095, 0),
		(drawing, 360, 360, 4095, 4095, 0),
		(drawing, 361, 361, 4095, 4095, 0),
		(drawing, 362, 362, 4095, 4095, 0),
		(drawing, 363, 363, 4095, 4095, 0),
		(drawing, 364, 364, 4095, 4095, 0),
		(drawing, 365, 365, 4095, 4095, 0),
		(drawing, 366, 366, 4095, 4095, 0),
		(drawing, 367, 367, 4095, 4095, 0),
		(drawing, 368, 368, 4095, 4095, 0),
		(drawing, 369, 369, 4095, 4095, 0),
		(drawing, 370, 370, 4095, 4095, 0),
		(drawing, 371, 371, 4095, 4095, 0),
		(drawing, 372, 372, 4095, 4095, 0),
		(drawing, 373, 373, 4095, 4095, 0),
		(drawing, 374, 374, 4095, 4095, 0),
		(drawing, 375, 375, 4095, 4095, 0),
		(drawing, 376, 376, 4095, 4095, 0),
		(drawing, 377, 377, 4095, 4095, 0),
		(drawing, 378, 378, 4095, 4095, 0),
		(drawing, 379, 379, 4095, 4095, 0),
		(drawing, 380, 380, 4095, 4095, 0),
		(drawing, 381, 381, 4095, 4095, 0),
		(drawing, 382, 382, 4095, 4095, 0),
		(drawing, 383, 383, 4095, 4095, 0),
		(drawing, 384, 384, 4095, 4095, 0),
		(drawing, 385, 385, 4095, 4095, 0),
		(drawing, 386, 386, 4095, 4095, 0),
		(drawing, 387, 387, 4095, 4095, 0),
		(drawing, 388, 388, 4095, 4095, 0),
		(drawing, 389, 389, 4095, 4095, 0),
		(drawing, 390, 390, 4095, 4095, 0),
		(drawing, 391, 391, 4095, 4095, 0),
		(drawing, 392, 392, 4095, 4095, 0),
		(drawing, 393, 393, 4095, 4095, 0),
		(drawing, 394, 394, 4095, 4095, 0),
		(drawing, 395, 395, 4095, 4095, 0),
		(drawing, 396, 396, 4095, 4095, 0),
		(drawing, 397, 397, 4095, 4095, 0),
		(drawing, 398, 398, 4095, 4095, 0),
		(drawing, 399, 399, 4095, 4095, 0),
		(drawing, 400, 400, 4095, 4095, 0),
		(drawing, 401, 401, 4095, 4095, 0),
		(drawing, 402, 402, 4095, 4095, 0),
		(drawing, 403, 403, 4095, 4095, 0),
		(drawing, 404, 404, 4095, 4095, 0),
		(drawing, 405, 405, 4095, 4095, 0),
		(drawing, 406, 406, 4095, 4095, 0),
		(drawing, 407, 407, 4095, 4095, 0),
		(drawing, 408, 408, 4095, 4095, 0),
		(drawing, 409, 409, 4095, 4095, 0),
		(drawing, 410, 410, 4095, 4095, 0),
		(drawing, 411, 411, 4095, 4095, 0),
		(drawing, 412, 412, 4095, 4095, 0),
		(drawing, 413, 413, 4095, 4095, 0),
		(drawing, 414, 414, 4095, 4095, 0),
		(drawing, 415, 415, 4095, 4095, 0),
		(drawing, 416, 416, 4095, 4095, 0),
		(drawing, 417, 417, 4095, 4095, 0),
		(drawing, 418, 418, 4095, 4095, 0),
		(drawing, 419, 419, 4095, 4095, 0),
		(drawing, 420, 420, 4095, 4095, 0),
		(drawing, 421, 421, 4095, 4095, 0),
		(drawing, 422, 422, 4095, 4095, 0),
		(drawing, 423, 423, 4095, 4095, 0),
		(drawing, 424, 424, 4095, 4095, 0),
		(drawing, 425, 425, 4095, 4095, 0),
		(drawing, 426, 426, 4095, 4095, 0),
		(drawing, 427, 427, 4095, 4095, 0),
		(drawing, 428, 428, 4095, 4095, 0),
		(drawing, 429, 429, 4095, 4095, 0),
		(drawing, 430, 430, 4095, 4095, 0),
		(drawing, 431, 431, 4095, 4095, 0),
		(drawing, 432, 432, 4095, 4095, 0),
		(drawing, 433, 433, 4095, 4095, 0),
		(drawing, 434, 434, 4095, 4095, 0),
		(drawing, 435, 435, 4095, 4095, 0),
		(drawing, 436, 436, 4095, 4095, 0),
		(drawing, 437, 437, 4095, 4095, 0),
		(drawing, 438, 438, 4095, 4095, 0),
		(drawing, 439, 439, 4095, 4095, 0),
		(drawing, 440, 440, 4095, 4095, 0),
		(drawing, 441, 441, 4095, 4095, 0),
		(drawing, 442, 442, 4095, 4095, 0),
		(drawing, 443, 443, 4095, 4095, 0),
		(drawing, 444, 444, 4095, 4095, 0),
		(drawing, 445, 445, 4095, 4095, 0),
		(drawing, 446, 446, 4095, 4095, 0),
		(drawing, 447, 447, 4095, 4095, 0),
		(drawing, 448, 448, 4095, 4095, 0),
		(drawing, 449, 449, 4095, 4095, 0),
		(drawing, 450, 450, 4095, 4095, 0),
		(drawing, 451, 451, 4095, 4095, 0),
		(drawing, 452, 452, 4095, 4095, 0),
		(drawing, 453, 453, 4095, 4095, 0),
		(drawing, 454, 454, 4095, 4095, 0),
		(drawing, 455, 455, 4095, 4095, 0),
		(drawing, 456, 456, 4095, 4095, 0),
		(drawing, 457, 457, 4095, 4095, 0),
		(drawing, 458, 458, 4095, 4095, 0),
		(drawing, 459, 459, 4095, 4095, 0),
		(drawing, 460, 460, 4095, 4095, 0),
		(drawing, 461, 461, 4095, 4095, 0),
		(drawing, 462, 462, 4095, 4095, 0),
		(drawing, 463, 463, 4095, 4095, 0),
		(drawing, 464, 464, 4095, 4095, 0),
		(drawing, 465, 465, 4095, 4095, 0),
		(drawing, 466, 466, 4095, 4095, 0),
		(drawing, 467, 467, 4095, 4095, 0),
		(drawing, 468, 468, 4095, 4095, 0),
		(drawing, 469, 469, 4095, 4095, 0),
		(drawing, 470, 470, 4095, 4095, 0),
		(drawing, 471, 471, 4095, 4095, 0),
		(drawing, 472, 472, 4095, 4095, 0),
		(drawing, 473, 473, 4095, 4095, 0),
		(drawing, 474, 474, 4095, 4095, 0),
		(drawing, 475, 475, 4095, 4095, 0),
		(drawing, 476, 476, 4095, 4095, 0),
		(drawing, 477, 477, 4095, 4095, 0),
		(drawing, 478, 478, 4095, 4095, 0),
		(drawing, 479, 479, 4095, 4095, 0),
		(drawing, 480, 480, 4095, 4095, 0),
		(drawing, 481, 481, 4095, 4095, 0),
		(drawing, 482, 482, 4095, 4095, 0),
		(drawing, 483, 483, 4095, 4095, 0),
		(drawing, 484, 484, 4095, 4095, 0),
		(drawing, 485, 485, 4095, 4095, 0),
		(drawing, 486, 486, 4095, 4095, 0),
		(drawing, 487, 487, 4095, 4095, 0),
		(drawing, 488, 488, 4095, 4095, 0),
		(drawing, 489, 489, 4095, 4095, 0),
		(drawing, 490, 490, 4095, 4095, 0),
		(drawing, 491, 491, 4095, 4095, 0),
		(drawing, 492, 492, 4095, 4095, 0),
		(drawing, 493, 493, 4095, 4095, 0),
		(drawing, 494, 494, 4095, 4095, 0),
		(drawing, 495, 495, 4095, 4095, 0),
		(drawing, 496, 496, 4095, 4095, 0),
		(drawing, 497, 497, 4095, 4095, 0),
		(drawing, 498, 498, 4095, 4095, 0),
		(drawing, 499, 499, 4095, 4095, 0),
		(drawing, 500, 500, 4095, 4095, 0),
		(drawing, 501, 501, 4095, 4095, 0),
		(drawing, 502, 502, 4095, 4095, 0),
		(drawing, 503, 503, 4095, 4095, 0),
		(drawing, 504, 504, 4095, 4095, 0),
		(drawing, 505, 505, 4095, 4095, 0),
		(drawing, 506, 506, 4095, 4095, 0),
		(drawing, 507, 507, 4095, 4095, 0),
		(drawing, 508, 508, 4095, 4095, 0),
		(drawing, 509, 509, 4095, 4095, 0),
		(drawing, 510, 510, 4095, 4095, 0),
		(drawing, 511, 511, 4095, 4095, 0),
		(drawing, 512, 512, 4095, 4095, 0),
		(drawing, 513, 513, 4095, 4095, 0),
		(drawing, 514, 514, 4095, 4095, 0),
		(drawing, 515, 515, 4095, 4095, 0),
		(drawing, 516, 516, 4095, 4095, 0),
		(drawing, 517, 517, 4095, 4095, 0),
		(drawing, 518, 518, 4095, 4095, 0),
		(drawing, 519, 519, 4095, 4095, 0),
		(drawing, 520, 520, 4095, 4095, 0),
		(drawing, 521, 521, 4095, 4095, 0),
		(drawing, 522, 522, 4095, 4095, 0),
		(drawing, 523, 523, 4095, 4095, 0),
		(drawing, 524, 524, 4095, 4095, 0),
		(drawing, 525, 525, 4095, 4095, 0),
		(drawing, 526, 526, 4095, 4095, 0),
		(drawing, 527, 527, 4095, 4095, 0),
		(drawing, 528, 528, 4095, 4095, 0),
		(drawing, 529, 529, 4095, 4095, 0),
		(drawing, 530, 530, 4095, 4095, 0),
		(drawing, 531, 531, 4095, 4095, 0),
		(drawing, 532, 532, 4095, 4095, 0),
		(drawing, 533, 533, 4095, 4095, 0),
		(drawing, 534, 534, 4095, 4095, 0),
		(drawing, 535, 535, 4095, 4095, 0),
		(drawing, 536, 536, 4095, 4095, 0),
		(drawing, 537, 537, 4095, 4095, 0),
		(drawing, 538, 538, 4095, 4095, 0),
		(drawing, 539, 539, 4095, 4095, 0),
		(drawing, 540, 540, 4095, 4095, 0),
		(drawing, 541, 541, 4095, 4095, 0),
		(drawing, 542, 542, 4095, 4095, 0),
		(drawing, 543, 543, 4095, 4095, 0),
		(drawing, 544, 544, 4095, 4095, 0),
		(drawing, 545, 545, 4095, 4095, 0),
		(drawing, 546, 546, 4095, 4095, 0),
		(drawing, 547, 547, 4095, 4095, 0),
		(drawing, 548, 548, 4095, 4095, 0),
		(drawing, 549, 549, 4095, 4095, 0),
		(drawing, 550, 550, 4095, 4095, 0),
		(drawing, 551, 551, 4095, 4095, 0),
		(drawing, 552, 552, 4095, 4095, 0),
		(drawing, 553, 553, 4095, 4095, 0),
		(drawing, 554, 554, 4095, 4095, 0),
		(drawing, 555, 555, 4095, 4095, 0),
		(drawing, 556, 556, 4095, 4095, 0),
		(drawing, 557, 557, 4095, 4095, 0),
		(drawing, 558, 558, 4095, 4095, 0),
		(drawing, 559, 559, 4095, 4095, 0),
		(drawing, 560, 560, 4095, 4095, 0),
		(drawing, 561, 561, 4095, 4095, 0),
		(drawing, 562, 562, 4095, 4095, 0),
		(drawing, 563, 563, 4095, 4095, 0),
		(drawing, 564, 564, 4095, 4095, 0),
		(drawing, 565, 565, 4095, 4095, 0),
		(drawing, 566, 566, 4095, 4095, 0),
		(drawing, 567, 567, 4095, 4095, 0),
		(drawing, 568, 568, 4095, 4095, 0),
		(drawing, 569, 569, 4095, 4095, 0),
		(drawing, 570, 570, 4095, 4095, 0),
		(drawing, 571, 571, 4095, 4095, 0),
		(drawing, 572, 572, 4095, 4095, 0),
		(drawing, 573, 573, 4095, 4095, 0),
		(drawing, 574, 574, 4095, 4095, 0),
		(drawing, 575, 575, 4095, 4095, 0),
		(drawing, 576, 576, 4095, 4095, 0),
		(drawing, 577, 577, 4095, 4095, 0),
		(drawing, 578, 578, 4095, 4095, 0),
		(drawing, 579, 579, 4095, 4095, 0),
		(drawing, 580, 580, 4095, 4095, 0),
		(drawing, 581, 581, 4095, 4095, 0),
		(drawing, 582, 582, 4095, 4095, 0),
		(drawing, 583, 583, 4095, 4095, 0),
		(drawing, 584, 584, 4095, 4095, 0),
		(drawing, 585, 585, 4095, 4095, 0),
		(drawing, 586, 586, 4095, 4095, 0),
		(drawing, 587, 587, 4095, 4095, 0),
		(drawing, 588, 588, 4095, 4095, 0),
		(drawing, 589, 589, 4095, 4095, 0),
		(drawing, 590, 590, 4095, 4095, 0),
		(drawing, 591, 591, 4095, 4095, 0),
		(drawing, 592, 592, 4095, 4095, 0),
		(drawing, 593, 593, 4095, 4095, 0),
		(drawing, 594, 594, 4095, 4095, 0),
		(drawing, 595, 595, 4095, 4095, 0),
		(drawing, 596, 596, 4095, 4095, 0),
		(drawing, 597, 597, 4095, 4095, 0),
		(drawing, 598, 598, 4095, 4095, 0),
		(drawing, 599, 599, 4095, 4095, 0),
		(drawing, 600, 600, 4095, 4095, 0),
		(drawing, 601, 601, 4095, 4095, 0),
		(drawing, 602, 602, 4095, 4095, 0),
		(drawing, 603, 603, 4095, 4095, 0),
		(drawing, 604, 604, 4095, 4095, 0),
		(drawing, 605, 605, 4095, 4095, 0),
		(drawing, 606, 606, 4095, 4095, 0),
		(drawing, 607, 607, 4095, 4095, 0),
		(drawing, 608, 608, 4095, 4095, 0),
		(drawing, 609, 609, 4095, 4095, 0),
		(drawing, 610, 610, 4095, 4095, 0),
		(drawing, 611, 611, 4095, 4095, 0),
		(drawing, 612, 612, 4095, 4095, 0),
		(drawing, 613, 613, 4095, 4095, 0),
		(drawing, 614, 614, 4095, 4095, 0),
		(drawing, 615, 615, 4095, 4095, 0),
		(drawing, 616, 616, 4095, 4095, 0),
		(drawing, 617, 617, 4095, 4095, 0),
		(drawing, 618, 618, 4095, 4095, 0),
		(drawing, 619, 619, 4095, 4095, 0),
		(drawing, 620, 620, 4095, 4095, 0),
		(drawing, 621, 621, 4095, 4095, 0),
		(drawing, 622, 622, 4095, 4095, 0),
		(drawing, 623, 623, 4095, 4095, 0),
		(drawing, 624, 624, 4095, 4095, 0),
		(drawing, 625, 625, 4095, 4095, 0),
		(drawing, 626, 626, 4095, 4095, 0),
		(drawing, 627, 627, 4095, 4095, 0),
		(drawing, 628, 628, 4095, 4095, 0),
		(drawing, 629, 629, 4095, 4095, 0),
		(drawing, 630, 630, 4095, 4095, 0),
		(drawing, 631, 631, 4095, 4095, 0),
		(drawing, 632, 632, 4095, 4095, 0),
		(drawing, 633, 633, 4095, 4095, 0),
		(drawing, 634, 634, 4095, 4095, 0),
		(drawing, 635, 635, 4095, 4095, 0),
		(drawing, 636, 636, 4095, 4095, 0),
		(drawing, 637, 637, 4095, 4095, 0),
		(drawing, 638, 638, 4095, 4095, 0),
		(drawing, 639, 639, 4095, 4095, 0),
		(drawing, 640, 640, 4095, 4095, 0),
		(drawing, 641, 641, 4095, 4095, 0),
		(drawing, 642, 642, 4095, 4095, 0),
		(drawing, 643, 643, 4095, 4095, 0),
		(drawing, 644, 644, 4095, 4095, 0),
		(drawing, 645, 645, 4095, 4095, 0),
		(drawing, 646, 646, 4095, 4095, 0),
		(drawing, 647, 647, 4095, 4095, 0),
		(drawing, 648, 648, 4095, 4095, 0),
		(drawing, 649, 649, 4095, 4095, 0),
		(drawing, 650, 650, 4095, 4095, 0),
		(drawing, 651, 651, 4095, 4095, 0),
		(drawing, 652, 652, 4095, 4095, 0),
		(drawing, 653, 653, 4095, 4095, 0),
		(drawing, 654, 654, 4095, 4095, 0),
		(drawing, 655, 655, 4095, 4095, 0),
		(drawing, 656, 656, 4095, 4095, 0),
		(drawing, 657, 657, 4095, 4095, 0),
		(drawing, 658, 658, 4095, 4095, 0),
		(drawing, 659, 659, 4095, 4095, 0),
		(drawing, 660, 660, 4095, 4095, 0),
		(drawing, 661, 661, 4095, 4095, 0),
		(drawing, 662, 662, 4095, 4095, 0),
		(drawing, 663, 663, 4095, 4095, 0),
		(drawing, 664, 664, 4095, 4095, 0),
		(drawing, 665, 665, 4095, 4095, 0),
		(drawing, 666, 666, 4095, 4095, 0),
		(drawing, 667, 667, 4095, 4095, 0),
		(drawing, 668, 668, 4095, 4095, 0),
		(drawing, 669, 669, 4095, 4095, 0),
		(drawing, 670, 670, 4095, 4095, 0),
		(drawing, 671, 671, 4095, 4095, 0),
		(drawing, 672, 672, 4095, 4095, 0),
		(drawing, 673, 673, 4095, 4095, 0),
		(drawing, 674, 674, 4095, 4095, 0),
		(drawing, 675, 675, 4095, 4095, 0),
		(drawing, 676, 676, 4095, 4095, 0),
		(drawing, 677, 677, 4095, 4095, 0),
		(drawing, 678, 678, 4095, 4095, 0),
		(drawing, 679, 679, 4095, 4095, 0),
		(drawing, 680, 680, 4095, 4095, 0),
		(drawing, 681, 681, 4095, 4095, 0),
		(drawing, 682, 682, 4095, 4095, 0),
		(drawing, 683, 683, 4095, 4095, 0),
		(drawing, 684, 684, 4095, 4095, 0),
		(drawing, 685, 685, 4095, 4095, 0),
		(drawing, 686, 686, 4095, 4095, 0),
		(drawing, 687, 687, 4095, 4095, 0),
		(drawing, 688, 688, 4095, 4095, 0),
		(drawing, 689, 689, 4095, 4095, 0),
		(drawing, 690, 690, 4095, 4095, 0),
		(drawing, 691, 691, 4095, 4095, 0),
		(drawing, 692, 692, 4095, 4095, 0),
		(drawing, 693, 693, 4095, 4095, 0),
		(drawing, 694, 694, 4095, 4095, 0),
		(drawing, 695, 695, 4095, 4095, 0),
		(drawing, 696, 696, 4095, 4095, 0),
		(drawing, 697, 697, 4095, 4095, 0),
		(drawing, 698, 698, 4095, 4095, 0),
		(drawing, 699, 699, 4095, 4095, 0),
		(drawing, 700, 700, 4095, 4095, 0),
		(drawing, 701, 701, 4095, 4095, 0),
		(drawing, 702, 702, 4095, 4095, 0),
		(drawing, 703, 703, 4095, 4095, 0),
		(drawing, 704, 704, 4095, 4095, 0),
		(drawing, 705, 705, 4095, 4095, 0),
		(drawing, 706, 706, 4095, 4095, 0),
		(drawing, 707, 707, 4095, 4095, 0),
		(drawing, 708, 708, 4095, 4095, 0),
		(drawing, 709, 709, 4095, 4095, 0),
		(drawing, 710, 710, 4095, 4095, 0),
		(drawing, 711, 711, 4095, 4095, 0),
		(drawing, 712, 712, 4095, 4095, 0),
		(drawing, 713, 713, 4095, 4095, 0),
		(drawing, 714, 714, 4095, 4095, 0),
		(drawing, 715, 715, 4095, 4095, 0),
		(drawing, 716, 716, 4095, 4095, 0),
		(drawing, 717, 717, 4095, 4095, 0),
		(drawing, 718, 718, 4095, 4095, 0),
		(drawing, 719, 719, 4095, 4095, 0),
		(drawing, 720, 720, 4095, 4095, 0),
		(drawing, 721, 721, 4095, 4095, 0),
		(drawing, 722, 722, 4095, 4095, 0),
		(drawing, 723, 723, 4095, 4095, 0),
		(drawing, 724, 724, 4095, 4095, 0),
		(drawing, 725, 725, 4095, 4095, 0),
		(drawing, 726, 726, 4095, 4095, 0),
		(drawing, 727, 727, 4095, 4095, 0),
		(drawing, 728, 728, 4095, 4095, 0),
		(drawing, 729, 729, 4095, 4095, 0),
		(drawing, 730, 730, 4095, 4095, 0),
		(drawing, 731, 731, 4095, 4095, 0),
		(drawing, 732, 732, 4095, 4095, 0),
		(drawing, 733, 733, 4095, 4095, 0),
		(drawing, 734, 734, 4095, 4095, 0),
		(drawing, 735, 735, 4095, 4095, 0),
		(drawing, 736, 736, 4095, 4095, 0),
		(drawing, 737, 737, 4095, 4095, 0),
		(drawing, 738, 738, 4095, 4095, 0),
		(drawing, 739, 739, 4095, 4095, 0),
		(drawing, 740, 740, 4095, 4095, 0),
		(drawing, 741, 741, 4095, 4095, 0),
		(drawing, 742, 742, 4095, 4095, 0),
		(drawing, 743, 743, 4095, 4095, 0),
		(drawing, 744, 744, 4095, 4095, 0),
		(drawing, 745, 745, 4095, 4095, 0),
		(drawing, 746, 746, 4095, 4095, 0),
		(drawing, 747, 747, 4095, 4095, 0),
		(drawing, 748, 748, 4095, 4095, 0),
		(drawing, 749, 749, 4095, 4095, 0),
		(drawing, 750, 750, 4095, 4095, 0),
		(drawing, 751, 751, 4095, 4095, 0),
		(drawing, 752, 752, 4095, 4095, 0),
		(drawing, 753, 753, 4095, 4095, 0),
		(drawing, 754, 754, 4095, 4095, 0),
		(drawing, 755, 755, 4095, 4095, 0),
		(drawing, 756, 756, 4095, 4095, 0),
		(drawing, 757, 757, 4095, 4095, 0),
		(drawing, 758, 758, 4095, 4095, 0),
		(drawing, 759, 759, 4095, 4095, 0),
		(drawing, 760, 760, 4095, 4095, 0),
		(drawing, 761, 761, 4095, 4095, 0),
		(drawing, 762, 762, 4095, 4095, 0),
		(drawing, 763, 763, 4095, 4095, 0),
		(drawing, 764, 764, 4095, 4095, 0),
		(drawing, 765, 765, 4095, 4095, 0),
		(drawing, 766, 766, 4095, 4095, 0),
		(drawing, 767, 767, 4095, 4095, 0),
		(drawing, 768, 768, 4095, 4095, 0),
		(drawing, 769, 769, 4095, 4095, 0),
		(drawing, 770, 770, 4095, 4095, 0),
		(drawing, 771, 771, 4095, 4095, 0),
		(drawing, 772, 772, 4095, 4095, 0),
		(drawing, 773, 773, 4095, 4095, 0),
		(drawing, 774, 774, 4095, 4095, 0),
		(drawing, 775, 775, 4095, 4095, 0),
		(drawing, 776, 776, 4095, 4095, 0),
		(drawing, 777, 777, 4095, 4095, 0),
		(drawing, 778, 778, 4095, 4095, 0),
		(drawing, 779, 779, 4095, 4095, 0),
		(drawing, 780, 780, 4095, 4095, 0),
		(drawing, 781, 781, 4095, 4095, 0),
		(drawing, 782, 782, 4095, 4095, 0),
		(drawing, 783, 783, 4095, 4095, 0),
		(drawing, 784, 784, 4095, 4095, 0),
		(drawing, 785, 785, 4095, 4095, 0),
		(drawing, 786, 786, 4095, 4095, 0),
		(drawing, 787, 787, 4095, 4095, 0),
		(drawing, 788, 788, 4095, 4095, 0),
		(drawing, 789, 789, 4095, 4095, 0),
		(drawing, 790, 790, 4095, 4095, 0),
		(drawing, 791, 791, 4095, 4095, 0),
		(drawing, 792, 792, 4095, 4095, 0),
		(drawing, 793, 793, 4095, 4095, 0),
		(drawing, 794, 794, 4095, 4095, 0),
		(drawing, 795, 795, 4095, 4095, 0),
		(drawing, 796, 796, 4095, 4095, 0),
		(drawing, 797, 797, 4095, 4095, 0),
		(drawing, 798, 798, 4095, 4095, 0),
		(drawing, 799, 799, 4095, 4095, 0),
		(drawing, 800, 800, 4095, 4095, 0),
		(drawing, 801, 801, 4095, 4095, 0),
		(drawing, 802, 802, 4095, 4095, 0),
		(drawing, 803, 803, 4095, 4095, 0),
		(drawing, 804, 804, 4095, 4095, 0),
		(drawing, 805, 805, 4095, 4095, 0),
		(drawing, 806, 806, 4095, 4095, 0),
		(drawing, 807, 807, 4095, 4095, 0),
		(drawing, 808, 808, 4095, 4095, 0),
		(drawing, 809, 809, 4095, 4095, 0),
		(drawing, 810, 810, 4095, 4095, 0),
		(drawing, 811, 811, 4095, 4095, 0),
		(drawing, 812, 812, 4095, 4095, 0),
		(drawing, 813, 813, 4095, 4095, 0),
		(drawing, 814, 814, 4095, 4095, 0),
		(drawing, 815, 815, 4095, 4095, 0),
		(drawing, 816, 816, 4095, 4095, 0),
		(drawing, 817, 817, 4095, 4095, 0),
		(drawing, 818, 818, 4095, 4095, 0),
		(drawing, 819, 819, 4095, 4095, 0),
		(drawing, 820, 820, 4095, 4095, 0),
		(drawing, 821, 821, 4095, 4095, 0),
		(drawing, 822, 822, 4095, 4095, 0),
		(drawing, 823, 823, 4095, 4095, 0),
		(drawing, 824, 824, 4095, 4095, 0),
		(drawing, 825, 825, 4095, 4095, 0),
		(drawing, 826, 826, 4095, 4095, 0),
		(drawing, 827, 827, 4095, 4095, 0),
		(drawing, 828, 828, 4095, 4095, 0),
		(drawing, 829, 829, 4095, 4095, 0),
		(drawing, 830, 830, 4095, 4095, 0),
		(drawing, 831, 831, 4095, 4095, 0),
		(drawing, 832, 832, 4095, 4095, 0),
		(drawing, 833, 833, 4095, 4095, 0),
		(drawing, 834, 834, 4095, 4095, 0),
		(drawing, 835, 835, 4095, 4095, 0),
		(drawing, 836, 836, 4095, 4095, 0),
		(drawing, 837, 837, 4095, 4095, 0),
		(drawing, 838, 838, 4095, 4095, 0),
		(drawing, 839, 839, 4095, 4095, 0),
		(drawing, 840, 840, 4095, 4095, 0),
		(drawing, 841, 841, 4095, 4095, 0),
		(drawing, 842, 842, 4095, 4095, 0),
		(drawing, 843, 843, 4095, 4095, 0),
		(drawing, 844, 844, 4095, 4095, 0),
		(drawing, 845, 845, 4095, 4095, 0),
		(drawing, 846, 846, 4095, 4095, 0),
		(drawing, 847, 847, 4095, 4095, 0),
		(drawing, 848, 848, 4095, 4095, 0),
		(drawing, 849, 849, 4095, 4095, 0),
		(drawing, 850, 850, 4095, 4095, 0),
		(drawing, 851, 851, 4095, 4095, 0),
		(drawing, 852, 852, 4095, 4095, 0),
		(drawing, 853, 853, 4095, 4095, 0),
		(drawing, 854, 854, 4095, 4095, 0),
		(drawing, 855, 855, 4095, 4095, 0),
		(drawing, 856, 856, 4095, 4095, 0),
		(drawing, 857, 857, 4095, 4095, 0),
		(drawing, 858, 858, 4095, 4095, 0),
		(drawing, 859, 859, 4095, 4095, 0),
		(drawing, 860, 860, 4095, 4095, 0),
		(drawing, 861, 861, 4095, 4095, 0),
		(drawing, 862, 862, 4095, 4095, 0),
		(drawing, 863, 863, 4095, 4095, 0),
		(drawing, 864, 864, 4095, 4095, 0),
		(drawing, 865, 865, 4095, 4095, 0),
		(drawing, 866, 866, 4095, 4095, 0),
		(drawing, 867, 867, 4095, 4095, 0),
		(drawing, 868, 868, 4095, 4095, 0),
		(drawing, 869, 869, 4095, 4095, 0),
		(drawing, 870, 870, 4095, 4095, 0),
		(drawing, 871, 871, 4095, 4095, 0),
		(drawing, 872, 872, 4095, 4095, 0),
		(drawing, 873, 873, 4095, 4095, 0),
		(drawing, 874, 874, 4095, 4095, 0),
		(drawing, 875, 875, 4095, 4095, 0),
		(drawing, 876, 876, 4095, 4095, 0),
		(drawing, 877, 877, 4095, 4095, 0),
		(drawing, 878, 878, 4095, 4095, 0),
		(drawing, 879, 879, 4095, 4095, 0),
		(drawing, 880, 880, 4095, 4095, 0),
		(drawing, 881, 881, 4095, 4095, 0),
		(drawing, 882, 882, 4095, 4095, 0),
		(drawing, 883, 883, 4095, 4095, 0),
		(drawing, 884, 884, 4095, 4095, 0),
		(drawing, 885, 885, 4095, 4095, 0),
		(drawing, 886, 886, 4095, 4095, 0),
		(drawing, 887, 887, 4095, 4095, 0),
		(drawing, 888, 888, 4095, 4095, 0),
		(drawing, 889, 889, 4095, 4095, 0),
		(drawing, 890, 890, 4095, 4095, 0),
		(drawing, 891, 891, 4095, 4095, 0),
		(drawing, 892, 892, 4095, 4095, 0),
		(drawing, 893, 893, 4095, 4095, 0),
		(drawing, 894, 894, 4095, 4095, 0),
		(drawing, 895, 895, 4095, 4095, 0),
		(drawing, 896, 896, 4095, 4095, 0),
		(drawing, 897, 897, 4095, 4095, 0),
		(drawing, 898, 898, 4095, 4095, 0),
		(drawing, 899, 899, 4095, 4095, 0),
		(drawing, 900, 900, 4095, 4095, 0),
		(drawing, 901, 901, 4095, 4095, 0),
		(drawing, 902, 902, 4095, 4095, 0),
		(drawing, 903, 903, 4095, 4095, 0),
		(drawing, 904, 904, 4095, 4095, 0),
		(drawing, 905, 905, 4095, 4095, 0),
		(drawing, 906, 906, 4095, 4095, 0),
		(drawing, 907, 907, 4095, 4095, 0),
		(drawing, 908, 908, 4095, 4095, 0),
		(drawing, 909, 909, 4095, 4095, 0),
		(drawing, 910, 910, 4095, 4095, 0),
		(drawing, 911, 911, 4095, 4095, 0),
		(drawing, 912, 912, 4095, 4095, 0),
		(drawing, 913, 913, 4095, 4095, 0),
		(drawing, 914, 914, 4095, 4095, 0),
		(drawing, 915, 915, 4095, 4095, 0),
		(drawing, 916, 916, 4095, 4095, 0),
		(drawing, 917, 917, 4095, 4095, 0),
		(drawing, 918, 918, 4095, 4095, 0),
		(drawing, 919, 919, 4095, 4095, 0),
		(drawing, 920, 920, 4095, 4095, 0),
		(drawing, 921, 921, 4095, 4095, 0),
		(drawing, 922, 922, 4095, 4095, 0),
		(drawing, 923, 923, 4095, 4095, 0),
		(drawing, 924, 924, 4095, 4095, 0),
		(drawing, 925, 925, 4095, 4095, 0),
		(drawing, 926, 926, 4095, 4095, 0),
		(drawing, 927, 927, 4095, 4095, 0),
		(drawing, 928, 928, 4095, 4095, 0),
		(drawing, 929, 929, 4095, 4095, 0),
		(drawing, 930, 930, 4095, 4095, 0),
		(drawing, 931, 931, 4095, 4095, 0),
		(drawing, 932, 932, 4095, 4095, 0),
		(drawing, 933, 933, 4095, 4095, 0),
		(drawing, 934, 934, 4095, 4095, 0),
		(drawing, 935, 935, 4095, 4095, 0),
		(drawing, 936, 936, 4095, 4095, 0),
		(drawing, 937, 937, 4095, 4095, 0),
		(drawing, 938, 938, 4095, 4095, 0),
		(drawing, 939, 939, 4095, 4095, 0),
		(drawing, 940, 940, 4095, 4095, 0),
		(drawing, 941, 941, 4095, 4095, 0),
		(drawing, 942, 942, 4095, 4095, 0),
		(drawing, 943, 943, 4095, 4095, 0),
		(drawing, 944, 944, 4095, 4095, 0),
		(drawing, 945, 945, 4095, 4095, 0),
		(drawing, 946, 946, 4095, 4095, 0),
		(drawing, 947, 947, 4095, 4095, 0),
		(drawing, 948, 948, 4095, 4095, 0),
		(drawing, 949, 949, 4095, 4095, 0),
		(drawing, 950, 950, 4095, 4095, 0),
		(drawing, 951, 951, 4095, 4095, 0),
		(drawing, 952, 952, 4095, 4095, 0),
		(drawing, 953, 953, 4095, 4095, 0),
		(drawing, 954, 954, 4095, 4095, 0),
		(drawing, 955, 955, 4095, 4095, 0),
		(drawing, 956, 956, 4095, 4095, 0),
		(drawing, 957, 957, 4095, 4095, 0),
		(drawing, 958, 958, 4095, 4095, 0),
		(drawing, 959, 959, 4095, 4095, 0),
		(drawing, 960, 960, 4095, 4095, 0),
		(drawing, 961, 961, 4095, 4095, 0),
		(drawing, 962, 962, 4095, 4095, 0),
		(drawing, 963, 963, 4095, 4095, 0),
		(drawing, 964, 964, 4095, 4095, 0),
		(drawing, 965, 965, 4095, 4095, 0),
		(drawing, 966, 966, 4095, 4095, 0),
		(drawing, 967, 967, 4095, 4095, 0),
		(drawing, 968, 968, 4095, 4095, 0),
		(drawing, 969, 969, 4095, 4095, 0),
		(drawing, 970, 970, 4095, 4095, 0),
		(drawing, 971, 971, 4095, 4095, 0),
		(drawing, 972, 972, 4095, 4095, 0),
		(drawing, 973, 973, 4095, 4095, 0),
		(drawing, 974, 974, 4095, 4095, 0),
		(drawing, 975, 975, 4095, 4095, 0),
		(drawing, 976, 976, 4095, 4095, 0),
		(drawing, 977, 977, 4095, 4095, 0),
		(drawing, 978, 978, 4095, 4095, 0),
		(drawing, 979, 979, 4095, 4095, 0),
		(drawing, 980, 980, 4095, 4095, 0),
		(drawing, 981, 981, 4095, 4095, 0),
		(drawing, 982, 982, 4095, 4095, 0),
		(drawing, 983, 983, 4095, 4095, 0),
		(drawing, 984, 984, 4095, 4095, 0),
		(drawing, 985, 985, 4095, 4095, 0),
		(drawing, 986, 986, 4095, 4095, 0),
		(drawing, 987, 987, 4095, 4095, 0),
		(drawing, 988, 988, 4095, 4095, 0),
		(drawing, 989, 989, 4095, 4095, 0),
		(drawing, 990, 990, 4095, 4095, 0),
		(drawing, 991, 991, 4095, 4095, 0),
		(drawing, 992, 992, 4095, 4095, 0),
		(drawing, 993, 993, 4095, 4095, 0),
		(drawing, 994, 994, 4095, 4095, 0),
		(drawing, 995, 995, 4095, 4095, 0),
		(drawing, 996, 996, 4095, 4095, 0),
		(drawing, 997, 997, 4095, 4095, 0),
		(drawing, 998, 998, 4095, 4095, 0),
		(drawing, 999, 999, 4095, 4095, 0),
		(drawing, 1000, 1000, 4095, 4095, 0),
		(drawing, 1001, 1001, 4095, 4095, 0),
		(drawing, 1002, 1002, 4095, 4095, 0),
		(drawing, 1003, 1003, 4095, 4095, 0),
		(drawing, 1004, 1004, 4095, 4095, 0),
		(drawing, 1005, 1005, 4095, 4095, 0),
		(drawing, 1006, 1006, 4095, 4095, 0),
		(drawing, 1007, 1007, 4095, 4095, 0),
		(drawing, 1008, 1008, 4095, 4095, 0),
		(drawing, 1009, 1009, 4095, 4095, 0),
		(drawing, 1010, 1010, 4095, 4095, 0),
		(drawing, 1011, 1011, 4095, 4095, 0),
		(drawing, 1012, 1012, 4095, 4095, 0),
		(drawing, 1013, 1013, 4095, 4095, 0),
		(drawing, 1014, 1014, 4095, 4095, 0),
		(drawing, 1015, 1015, 4095, 4095, 0),
		(drawing, 1016, 1016, 4095, 4095, 0),
		(drawing, 1017, 1017, 4095, 4095, 0),
		(drawing, 1018, 1018, 4095, 4095, 0),
		(drawing, 1019, 1019, 4095, 4095, 0),
		(drawing, 1020, 1020, 4095, 4095, 0),
		(drawing, 1021, 1021, 4095, 4095, 0),
		(drawing, 1022, 1022, 4095, 4095, 0),
		(drawing, 1023, 1023, 4095, 4095, 0),
		(drawing, 1024, 1024, 4095, 4095, 0),
		(drawing, 1025, 1025, 4095, 4095, 0),
		(drawing, 1026, 1026, 4095, 4095, 0),
		(drawing, 1027, 1027, 4095, 4095, 0),
		(drawing, 1028, 1028, 4095, 4095, 0),
		(drawing, 1029, 1029, 4095, 4095, 0),
		(drawing, 1030, 1030, 4095, 4095, 0),
		(drawing, 1031, 1031, 4095, 4095, 0),
		(drawing, 1032, 1032, 4095, 4095, 0),
		(drawing, 1033, 1033, 4095, 4095, 0),
		(drawing, 1034, 1034, 4095, 4095, 0),
		(drawing, 1035, 1035, 4095, 4095, 0),
		(drawing, 1036, 1036, 4095, 4095, 0),
		(drawing, 1037, 1037, 4095, 4095, 0),
		(drawing, 1038, 1038, 4095, 4095, 0),
		(drawing, 1039, 1039, 4095, 4095, 0),
		(drawing, 1040, 1040, 4095, 4095, 0),
		(drawing, 1041, 1041, 4095, 4095, 0),
		(drawing, 1042, 1042, 4095, 4095, 0),
		(drawing, 1043, 1043, 4095, 4095, 0),
		(drawing, 1044, 1044, 4095, 4095, 0),
		(drawing, 1045, 1045, 4095, 4095, 0),
		(drawing, 1046, 1046, 4095, 4095, 0),
		(drawing, 1047, 1047, 4095, 4095, 0),
		(drawing, 1048, 1048, 4095, 4095, 0),
		(drawing, 1049, 1049, 4095, 4095, 0),
		(drawing, 1050, 1050, 4095, 4095, 0),
		(drawing, 1051, 1051, 4095, 4095, 0),
		(drawing, 1052, 1052, 4095, 4095, 0),
		(drawing, 1053, 1053, 4095, 4095, 0),
		(drawing, 1054, 1054, 4095, 4095, 0),
		(drawing, 1055, 1055, 4095, 4095, 0),
		(drawing, 1056, 1056, 4095, 4095, 0),
		(drawing, 1057, 1057, 4095, 4095, 0),
		(drawing, 1058, 1058, 4095, 4095, 0),
		(drawing, 1059, 1059, 4095, 4095, 0),
		(drawing, 1060, 1060, 4095, 4095, 0),
		(drawing, 1061, 1061, 4095, 4095, 0),
		(drawing, 1062, 1062, 4095, 4095, 0),
		(drawing, 1063, 1063, 4095, 4095, 0),
		(drawing, 1064, 1064, 4095, 4095, 0),
		(drawing, 1065, 1065, 4095, 4095, 0),
		(drawing, 1066, 1066, 4095, 4095, 0),
		(drawing, 1067, 1067, 4095, 4095, 0),
		(drawing, 1068, 1068, 4095, 4095, 0),
		(drawing, 1069, 1069, 4095, 4095, 0),
		(drawing, 1070, 1070, 4095, 4095, 0),
		(drawing, 1071, 1071, 4095, 4095, 0),
		(drawing, 1072, 1072, 4095, 4095, 0),
		(drawing, 1073, 1073, 4095, 4095, 0),
		(drawing, 1074, 1074, 4095, 4095, 0),
		(drawing, 1075, 1075, 4095, 4095, 0),
		(drawing, 1076, 1076, 4095, 4095, 0),
		(drawing, 1077, 1077, 4095, 4095, 0),
		(drawing, 1078, 1078, 4095, 4095, 0),
		(drawing, 1079, 1079, 4095, 4095, 0),
		(drawing, 1080, 1080, 4095, 4095, 0),
		(drawing, 1081, 1081, 4095, 4095, 0),
		(drawing, 1082, 1082, 4095, 4095, 0),
		(drawing, 1083, 1083, 4095, 4095, 0),
		(drawing, 1084, 1084, 4095, 4095, 0),
		(drawing, 1085, 1085, 4095, 4095, 0),
		(drawing, 1086, 1086, 4095, 4095, 0),
		(drawing, 1087, 1087, 4095, 4095, 0),
		(drawing, 1088, 1088, 4095, 4095, 0),
		(drawing, 1089, 1089, 4095, 4095, 0),
		(drawing, 1090, 1090, 4095, 4095, 0),
		(drawing, 1091, 1091, 4095, 4095, 0),
		(drawing, 1092, 1092, 4095, 4095, 0),
		(drawing, 1093, 1093, 4095, 4095, 0),
		(drawing, 1094, 1094, 4095, 4095, 0),
		(drawing, 1095, 1095, 4095, 4095, 0),
		(drawing, 1096, 1096, 4095, 4095, 0),
		(drawing, 1097, 1097, 4095, 4095, 0),
		(drawing, 1098, 1098, 4095, 4095, 0),
		(drawing, 1099, 1099, 4095, 4095, 0),
		(drawing, 1100, 1100, 4095, 4095, 0),
		(drawing, 1101, 1101, 4095, 4095, 0),
		(drawing, 1102, 1102, 4095, 4095, 0),
		(drawing, 1103, 1103, 4095, 4095, 0),
		(drawing, 1104, 1104, 4095, 4095, 0),
		(drawing, 1105, 1105, 4095, 4095, 0),
		(drawing, 1106, 1106, 4095, 4095, 0),
		(drawing, 1107, 1107, 4095, 4095, 0),
		(drawing, 1108, 1108, 4095, 4095, 0),
		(drawing, 1109, 1109, 4095, 4095, 0),
		(drawing, 1110, 1110, 4095, 4095, 0),
		(drawing, 1111, 1111, 4095, 4095, 0),
		(drawing, 1112, 1112, 4095, 4095, 0),
		(drawing, 1113, 1113, 4095, 4095, 0),
		(drawing, 1114, 1114, 4095, 4095, 0),
		(drawing, 1115, 1115, 4095, 4095, 0),
		(drawing, 1116, 1116, 4095, 4095, 0),
		(drawing, 1117, 1117, 4095, 4095, 0),
		(drawing, 1118, 1118, 4095, 4095, 0),
		(drawing, 1119, 1119, 4095, 4095, 0),
		(drawing, 1120, 1120, 4095, 4095, 0),
		(drawing, 1121, 1121, 4095, 4095, 0),
		(drawing, 1122, 1122, 4095, 4095, 0),
		(drawing, 1123, 1123, 4095, 4095, 0),
		(drawing, 1124, 1124, 4095, 4095, 0),
		(drawing, 1125, 1125, 4095, 4095, 0),
		(drawing, 1126, 1126, 4095, 4095, 0),
		(drawing, 1127, 1127, 4095, 4095, 0),
		(drawing, 1128, 1128, 4095, 4095, 0),
		(drawing, 1129, 1129, 4095, 4095, 0),
		(drawing, 1130, 1130, 4095, 4095, 0),
		(drawing, 1131, 1131, 4095, 4095, 0),
		(drawing, 1132, 1132, 4095, 4095, 0),
		(drawing, 1133, 1133, 4095, 4095, 0),
		(drawing, 1134, 1134, 4095, 4095, 0),
		(drawing, 1135, 1135, 4095, 4095, 0),
		(drawing, 1136, 1136, 4095, 4095, 0),
		(drawing, 1137, 1137, 4095, 4095, 0),
		(drawing, 1138, 1138, 4095, 4095, 0),
		(drawing, 1139, 1139, 4095, 4095, 0),
		(drawing, 1140, 1140, 4095, 4095, 0),
		(drawing, 1141, 1141, 4095, 4095, 0),
		(drawing, 1142, 1142, 4095, 4095, 0),
		(drawing, 1143, 1143, 4095, 4095, 0),
		(drawing, 1144, 1144, 4095, 4095, 0),
		(drawing, 1145, 1145, 4095, 4095, 0),
		(drawing, 1146, 1146, 4095, 4095, 0),
		(drawing, 1147, 1147, 4095, 4095, 0),
		(drawing, 1148, 1148, 4095, 4095, 0),
		(drawing, 1149, 1149, 4095, 4095, 0),
		(drawing, 1150, 1150, 4095, 4095, 0),
		(drawing, 1151, 1151, 4095, 4095, 0),
		(drawing, 1152, 1152, 4095, 4095, 0),
		(drawing, 1153, 1153, 4095, 4095, 0),
		(drawing, 1154, 1154, 4095, 4095, 0),
		(drawing, 1155, 1155, 4095, 4095, 0),
		(drawing, 1156, 1156, 4095, 4095, 0),
		(drawing, 1157, 1157, 4095, 4095, 0),
		(drawing, 1158, 1158, 4095, 4095, 0),
		(drawing, 1159, 1159, 4095, 4095, 0),
		(drawing, 1160, 1160, 4095, 4095, 0),
		(drawing, 1161, 1161, 4095, 4095, 0),
		(drawing, 1162, 1162, 4095, 4095, 0),
		(drawing, 1163, 1163, 4095, 4095, 0),
		(drawing, 1164, 1164, 4095, 4095, 0),
		(drawing, 1165, 1165, 4095, 4095, 0),
		(drawing, 1166, 1166, 4095, 4095, 0),
		(drawing, 1167, 1167, 4095, 4095, 0),
		(drawing, 1168, 1168, 4095, 4095, 0),
		(drawing, 1169, 1169, 4095, 4095, 0),
		(drawing, 1170, 1170, 4095, 4095, 0),
		(drawing, 1171, 1171, 4095, 4095, 0),
		(drawing, 1172, 1172, 4095, 4095, 0),
		(drawing, 1173, 1173, 4095, 4095, 0),
		(drawing, 1174, 1174, 4095, 4095, 0),
		(drawing, 1175, 1175, 4095, 4095, 0),
		(drawing, 1176, 1176, 4095, 4095, 0),
		(drawing, 1177, 1177, 4095, 4095, 0),
		(drawing, 1178, 1178, 4095, 4095, 0),
		(drawing, 1179, 1179, 4095, 4095, 0),
		(drawing, 1180, 1180, 4095, 4095, 0),
		(drawing, 1181, 1181, 4095, 4095, 0),
		(drawing, 1182, 1182, 4095, 4095, 0),
		(drawing, 1183, 1183, 4095, 4095, 0),
		(drawing, 1184, 1184, 4095, 4095, 0),
		(drawing, 1185, 1185, 4095, 4095, 0),
		(drawing, 1186, 1186, 4095, 4095, 0),
		(drawing, 1187, 1187, 4095, 4095, 0),
		(drawing, 1188, 1188, 4095, 4095, 0),
		(drawing, 1189, 1189, 4095, 4095, 0),
		(drawing, 1190, 1190, 4095, 4095, 0),
		(drawing, 1191, 1191, 4095, 4095, 0),
		(drawing, 1192, 1192, 4095, 4095, 0),
		(drawing, 1193, 1193, 4095, 4095, 0),
		(drawing, 1194, 1194, 4095, 4095, 0),
		(drawing, 1195, 1195, 4095, 4095, 0),
		(drawing, 1196, 1196, 4095, 4095, 0),
		(drawing, 1197, 1197, 4095, 4095, 0),
		(drawing, 1198, 1198, 4095, 4095, 0),
		(drawing, 1199, 1199, 4095, 4095, 0),
		(drawing, 1200, 1200, 4095, 4095, 0),
		(drawing, 1201, 1201, 4095, 4095, 0),
		(drawing, 1202, 1202, 4095, 4095, 0),
		(drawing, 1203, 1203, 4095, 4095, 0),
		(drawing, 1204, 1204, 4095, 4095, 0),
		(drawing, 1205, 1205, 4095, 4095, 0),
		(drawing, 1206, 1206, 4095, 4095, 0),
		(drawing, 1207, 1207, 4095, 4095, 0),
		(drawing, 1208, 1208, 4095, 4095, 0),
		(drawing, 1209, 1209, 4095, 4095, 0),
		(drawing, 1210, 1210, 4095, 4095, 0),
		(drawing, 1211, 1211, 4095, 4095, 0),
		(drawing, 1212, 1212, 4095, 4095, 0),
		(drawing, 1213, 1213, 4095, 4095, 0),
		(drawing, 1214, 1214, 4095, 4095, 0),
		(drawing, 1215, 1215, 4095, 4095, 0),
		(drawing, 1216, 1216, 4095, 4095, 0),
		(drawing, 1217, 1217, 4095, 4095, 0),
		(drawing, 1218, 1218, 4095, 4095, 0),
		(drawing, 1219, 1219, 4095, 4095, 0),
		(drawing, 1220, 1220, 4095, 4095, 0),
		(drawing, 1221, 1221, 4095, 4095, 0),
		(drawing, 1222, 1222, 4095, 4095, 0),
		(drawing, 1223, 1223, 4095, 4095, 0),
		(drawing, 1224, 1224, 4095, 4095, 0),
		(drawing, 1225, 1225, 4095, 4095, 0),
		(drawing, 1226, 1226, 4095, 4095, 0),
		(drawing, 1227, 1227, 4095, 4095, 0),
		(drawing, 1228, 1228, 4095, 4095, 0),
		(drawing, 1229, 1229, 4095, 4095, 0),
		(drawing, 1230, 1230, 4095, 4095, 0),
		(drawing, 1231, 1231, 4095, 4095, 0),
		(drawing, 1232, 1232, 4095, 4095, 0),
		(drawing, 1233, 1233, 4095, 4095, 0),
		(drawing, 1234, 1234, 4095, 4095, 0),
		(drawing, 1235, 1235, 4095, 4095, 0),
		(drawing, 1236, 1236, 4095, 4095, 0),
		(drawing, 1237, 1237, 4095, 4095, 0),
		(drawing, 1238, 1238, 4095, 4095, 0),
		(drawing, 1239, 1239, 4095, 4095, 0),
		(drawing, 1240, 1240, 4095, 4095, 0),
		(drawing, 1241, 1241, 4095, 4095, 0),
		(drawing, 1242, 1242, 4095, 4095, 0),
		(drawing, 1243, 1243, 4095, 4095, 0),
		(drawing, 1244, 1244, 4095, 4095, 0),
		(drawing, 1245, 1245, 4095, 4095, 0),
		(drawing, 1246, 1246, 4095, 4095, 0),
		(drawing, 1247, 1247, 4095, 4095, 0),
		(drawing, 1248, 1248, 4095, 4095, 0),
		(drawing, 1249, 1249, 4095, 4095, 0),
		(drawing, 1250, 1250, 4095, 4095, 0),
		(drawing, 1251, 1251, 4095, 4095, 0),
		(drawing, 1252, 1252, 4095, 4095, 0),
		(drawing, 1253, 1253, 4095, 4095, 0),
		(drawing, 1254, 1254, 4095, 4095, 0),
		(drawing, 1255, 1255, 4095, 4095, 0),
		(drawing, 1256, 1256, 4095, 4095, 0),
		(drawing, 1257, 1257, 4095, 4095, 0),
		(drawing, 1258, 1258, 4095, 4095, 0),
		(drawing, 1259, 1259, 4095, 4095, 0),
		(drawing, 1260, 1260, 4095, 4095, 0),
		(drawing, 1261, 1261, 4095, 4095, 0),
		(drawing, 1262, 1262, 4095, 4095, 0),
		(drawing, 1263, 1263, 4095, 4095, 0),
		(drawing, 1264, 1264, 4095, 4095, 0),
		(drawing, 1265, 1265, 4095, 4095, 0),
		(drawing, 1266, 1266, 4095, 4095, 0),
		(drawing, 1267, 1267, 4095, 4095, 0),
		(drawing, 1268, 1268, 4095, 4095, 0),
		(drawing, 1269, 1269, 4095, 4095, 0),
		(drawing, 1270, 1270, 4095, 4095, 0),
		(drawing, 1271, 1271, 4095, 4095, 0),
		(drawing, 1272, 1272, 4095, 4095, 0),
		(drawing, 1273, 1273, 4095, 4095, 0),
		(drawing, 1274, 1274, 4095, 4095, 0),
		(drawing, 1275, 1275, 4095, 4095, 0),
		(drawing, 1276, 1276, 4095, 4095, 0),
		(drawing, 1277, 1277, 4095, 4095, 0),
		(drawing, 1278, 1278, 4095, 4095, 0),
		(drawing, 1279, 1279, 4095, 4095, 0),
		(drawing, 1280, 1280, 4095, 4095, 0),
		(drawing, 1281, 1281, 4095, 4095, 0),
		(drawing, 1282, 1282, 4095, 4095, 0),
		(drawing, 1283, 1283, 4095, 4095, 0),
		(drawing, 1284, 1284, 4095, 4095, 0),
		(drawing, 1285, 1285, 4095, 4095, 0),
		(drawing, 1286, 1286, 4095, 4095, 0),
		(drawing, 1287, 1287, 4095, 4095, 0),
		(drawing, 1288, 1288, 4095, 4095, 0),
		(drawing, 1289, 1289, 4095, 4095, 0),
		(drawing, 1290, 1290, 4095, 4095, 0),
		(drawing, 1291, 1291, 4095, 4095, 0),
		(drawing, 1292, 1292, 4095, 4095, 0),
		(drawing, 1293, 1293, 4095, 4095, 0),
		(drawing, 1294, 1294, 4095, 4095, 0),
		(drawing, 1295, 1295, 4095, 4095, 0),
		(drawing, 1296, 1296, 4095, 4095, 0),
		(drawing, 1297, 1297, 4095, 4095, 0),
		(drawing, 1298, 1298, 4095, 4095, 0),
		(drawing, 1299, 1299, 4095, 4095, 0),
		(drawing, 1300, 1300, 4095, 4095, 0),
		(drawing, 1301, 1301, 4095, 4095, 0),
		(drawing, 1302, 1302, 4095, 4095, 0),
		(drawing, 1303, 1303, 4095, 4095, 0),
		(drawing, 1304, 1304, 4095, 4095, 0),
		(drawing, 1305, 1305, 4095, 4095, 0),
		(drawing, 1306, 1306, 4095, 4095, 0),
		(drawing, 1307, 1307, 4095, 4095, 0),
		(drawing, 1308, 1308, 4095, 4095, 0),
		(drawing, 1309, 1309, 4095, 4095, 0),
		(drawing, 1310, 1310, 4095, 4095, 0),
		(drawing, 1311, 1311, 4095, 4095, 0),
		(drawing, 1312, 1312, 4095, 4095, 0),
		(drawing, 1313, 1313, 4095, 4095, 0),
		(drawing, 1314, 1314, 4095, 4095, 0),
		(drawing, 1315, 1315, 4095, 4095, 0),
		(drawing, 1316, 1316, 4095, 4095, 0),
		(drawing, 1317, 1317, 4095, 4095, 0),
		(drawing, 1318, 1318, 4095, 4095, 0),
		(drawing, 1319, 1319, 4095, 4095, 0),
		(drawing, 1320, 1320, 4095, 4095, 0),
		(drawing, 1321, 1321, 4095, 4095, 0),
		(drawing, 1322, 1322, 4095, 4095, 0),
		(drawing, 1323, 1323, 4095, 4095, 0),
		(drawing, 1324, 1324, 4095, 4095, 0),
		(drawing, 1325, 1325, 4095, 4095, 0),
		(drawing, 1326, 1326, 4095, 4095, 0),
		(drawing, 1327, 1327, 4095, 4095, 0),
		(drawing, 1328, 1328, 4095, 4095, 0),
		(drawing, 1329, 1329, 4095, 4095, 0),
		(drawing, 1330, 1330, 4095, 4095, 0),
		(drawing, 1331, 1331, 4095, 4095, 0),
		(drawing, 1332, 1332, 4095, 4095, 0),
		(drawing, 1333, 1333, 4095, 4095, 0),
		(drawing, 1334, 1334, 4095, 4095, 0),
		(drawing, 1335, 1335, 4095, 4095, 0),
		(drawing, 1336, 1336, 4095, 4095, 0),
		(drawing, 1337, 1337, 4095, 4095, 0),
		(drawing, 1338, 1338, 4095, 4095, 0),
		(drawing, 1339, 1339, 4095, 4095, 0),
		(drawing, 1340, 1340, 4095, 4095, 0),
		(drawing, 1341, 1341, 4095, 4095, 0),
		(drawing, 1342, 1342, 4095, 4095, 0),
		(drawing, 1343, 1343, 4095, 4095, 0),
		(drawing, 1344, 1344, 4095, 4095, 0),
		(drawing, 1345, 1345, 4095, 4095, 0),
		(drawing, 1346, 1346, 4095, 4095, 0),
		(drawing, 1347, 1347, 4095, 4095, 0),
		(drawing, 1348, 1348, 4095, 4095, 0),
		(drawing, 1349, 1349, 4095, 4095, 0),
		(drawing, 1350, 1350, 4095, 4095, 0),
		(drawing, 1351, 1351, 4095, 4095, 0),
		(drawing, 1352, 1352, 4095, 4095, 0),
		(drawing, 1353, 1353, 4095, 4095, 0),
		(drawing, 1354, 1354, 4095, 4095, 0),
		(drawing, 1355, 1355, 4095, 4095, 0),
		(drawing, 1356, 1356, 4095, 4095, 0),
		(drawing, 1357, 1357, 4095, 4095, 0),
		(drawing, 1358, 1358, 4095, 4095, 0),
		(drawing, 1359, 1359, 4095, 4095, 0),
		(drawing, 1360, 1360, 4095, 4095, 0),
		(drawing, 1361, 1361, 4095, 4095, 0),
		(drawing, 1362, 1362, 4095, 4095, 0),
		(drawing, 1363, 1363, 4095, 4095, 0),
		(drawing, 1364, 1364, 4095, 4095, 0),
		(drawing, 1365, 1365, 4095, 4095, 0),
		(drawing, 1366, 1366, 4095, 4095, 0),
		(drawing, 1367, 1367, 4095, 4095, 0),
		(drawing, 1368, 1368, 4095, 4095, 0),
		(drawing, 1369, 1369, 4095, 4095, 0),
		(drawing, 1370, 1370, 4095, 4095, 0),
		(drawing, 1371, 1371, 4095, 4095, 0),
		(drawing, 1372, 1372, 4095, 4095, 0),
		(drawing, 1373, 1373, 4095, 4095, 0),
		(drawing, 1374, 1374, 4095, 4095, 0),
		(drawing, 1375, 1375, 4095, 4095, 0),
		(drawing, 1376, 1376, 4095, 4095, 0),
		(drawing, 1377, 1377, 4095, 4095, 0),
		(drawing, 1378, 1378, 4095, 4095, 0),
		(drawing, 1379, 1379, 4095, 4095, 0),
		(drawing, 1380, 1380, 4095, 4095, 0),
		(drawing, 1381, 1381, 4095, 4095, 0),
		(drawing, 1382, 1382, 4095, 4095, 0),
		(drawing, 1383, 1383, 4095, 4095, 0),
		(drawing, 1384, 1384, 4095, 4095, 0),
		(drawing, 1385, 1385, 4095, 4095, 0),
		(drawing, 1386, 1386, 4095, 4095, 0),
		(drawing, 1387, 1387, 4095, 4095, 0),
		(drawing, 1388, 1388, 4095, 4095, 0),
		(drawing, 1389, 1389, 4095, 4095, 0),
		(drawing, 1390, 1390, 4095, 4095, 0),
		(drawing, 1391, 1391, 4095, 4095, 0),
		(drawing, 1392, 1392, 4095, 4095, 0),
		(drawing, 1393, 1393, 4095, 4095, 0),
		(drawing, 1394, 1394, 4095, 4095, 0),
		(drawing, 1395, 1395, 4095, 4095, 0),
		(drawing, 1396, 1396, 4095, 4095, 0),
		(drawing, 1397, 1397, 4095, 4095, 0),
		(drawing, 1398, 1398, 4095, 4095, 0),
		(drawing, 1399, 1399, 4095, 4095, 0),
		(drawing, 1400, 1400, 4095, 4095, 0),
		(drawing, 1401, 1401, 4095, 4095, 0),
		(drawing, 1402, 1402, 4095, 4095, 0),
		(drawing, 1403, 1403, 4095, 4095, 0),
		(drawing, 1404, 1404, 4095, 4095, 0),
		(drawing, 1405, 1405, 4095, 4095, 0),
		(drawing, 1406, 1406, 4095, 4095, 0),
		(drawing, 1407, 1407, 4095, 4095, 0),
		(drawing, 1408, 1408, 4095, 4095, 0),
		(drawing, 1409, 1409, 4095, 4095, 0),
		(drawing, 1410, 1410, 4095, 4095, 0),
		(drawing, 1411, 1411, 4095, 4095, 0),
		(drawing, 1412, 1412, 4095, 4095, 0),
		(drawing, 1413, 1413, 4095, 4095, 0),
		(drawing, 1414, 1414, 4095, 4095, 0),
		(drawing, 1415, 1415, 4095, 4095, 0),
		(drawing, 1416, 1416, 4095, 4095, 0),
		(drawing, 1417, 1417, 4095, 4095, 0),
		(drawing, 1418, 1418, 4095, 4095, 0),
		(drawing, 1419, 1419, 4095, 4095, 0),
		(drawing, 1420, 1420, 4095, 4095, 0),
		(drawing, 1421, 1421, 4095, 4095, 0),
		(drawing, 1422, 1422, 4095, 4095, 0),
		(drawing, 1423, 1423, 4095, 4095, 0),
		(drawing, 1424, 1424, 4095, 4095, 0),
		(drawing, 1425, 1425, 4095, 4095, 0),
		(drawing, 1426, 1426, 4095, 4095, 0),
		(drawing, 1427, 1427, 4095, 4095, 0),
		(drawing, 1428, 1428, 4095, 4095, 0),
		(drawing, 1429, 1429, 4095, 4095, 0),
		(drawing, 1430, 1430, 4095, 4095, 0),
		(drawing, 1431, 1431, 4095, 4095, 0),
		(drawing, 1432, 1432, 4095, 4095, 0),
		(drawing, 1433, 1433, 4095, 4095, 0),
		(drawing, 1434, 1434, 4095, 4095, 0),
		(drawing, 1435, 1435, 4095, 4095, 0),
		(drawing, 1436, 1436, 4095, 4095, 0),
		(drawing, 1437, 1437, 4095, 4095, 0),
		(drawing, 1438, 1438, 4095, 4095, 0),
		(drawing, 1439, 1439, 4095, 4095, 0),
		(drawing, 1440, 1440, 4095, 4095, 0),
		(drawing, 1441, 1441, 4095, 4095, 0),
		(drawing, 1442, 1442, 4095, 4095, 0),
		(drawing, 1443, 1443, 4095, 4095, 0),
		(drawing, 1444, 1444, 4095, 4095, 0),
		(drawing, 1445, 1445, 4095, 4095, 0),
		(drawing, 1446, 1446, 4095, 4095, 0),
		(drawing, 1447, 1447, 4095, 4095, 0),
		(drawing, 1448, 1448, 4095, 4095, 0),
		(drawing, 1449, 1449, 4095, 4095, 0),
		(drawing, 1450, 1450, 4095, 4095, 0),
		(drawing, 1451, 1451, 4095, 4095, 0),
		(drawing, 1452, 1452, 4095, 4095, 0),
		(drawing, 1453, 1453, 4095, 4095, 0),
		(drawing, 1454, 1454, 4095, 4095, 0),
		(drawing, 1455, 1455, 4095, 4095, 0),
		(drawing, 1456, 1456, 4095, 4095, 0),
		(drawing, 1457, 1457, 4095, 4095, 0),
		(drawing, 1458, 1458, 4095, 4095, 0),
		(drawing, 1459, 1459, 4095, 4095, 0),
		(drawing, 1460, 1460, 4095, 4095, 0),
		(drawing, 1461, 1461, 4095, 4095, 0),
		(drawing, 1462, 1462, 4095, 4095, 0),
		(drawing, 1463, 1463, 4095, 4095, 0),
		(drawing, 1464, 1464, 4095, 4095, 0),
		(drawing, 1465, 1465, 4095, 4095, 0),
		(drawing, 1466, 1466, 4095, 4095, 0),
		(drawing, 1467, 1467, 4095, 4095, 0),
		(drawing, 1468, 1468, 4095, 4095, 0),
		(drawing, 1469, 1469, 4095, 4095, 0),
		(drawing, 1470, 1470, 4095, 4095, 0),
		(drawing, 1471, 1471, 4095, 4095, 0),
		(drawing, 1472, 1472, 4095, 4095, 0),
		(drawing, 1473, 1473, 4095, 4095, 0),
		(drawing, 1474, 1474, 4095, 4095, 0),
		(drawing, 1475, 1475, 4095, 4095, 0),
		(drawing, 1476, 1476, 4095, 4095, 0),
		(drawing, 1477, 1477, 4095, 4095, 0),
		(drawing, 1478, 1478, 4095, 4095, 0),
		(drawing, 1479, 1479, 4095, 4095, 0),
		(drawing, 1480, 1480, 4095, 4095, 0),
		(drawing, 1481, 1481, 4095, 4095, 0),
		(drawing, 1482, 1482, 4095, 4095, 0),
		(drawing, 1483, 1483, 4095, 4095, 0),
		(drawing, 1484, 1484, 4095, 4095, 0),
		(drawing, 1485, 1485, 4095, 4095, 0),
		(drawing, 1486, 1486, 4095, 4095, 0),
		(drawing, 1487, 1487, 4095, 4095, 0),
		(drawing, 1488, 1488, 4095, 4095, 0),
		(drawing, 1489, 1489, 4095, 4095, 0),
		(drawing, 1490, 1490, 4095, 4095, 0),
		(drawing, 1491, 1491, 4095, 4095, 0),
		(drawing, 1492, 1492, 4095, 4095, 0),
		(drawing, 1493, 1493, 4095, 4095, 0),
		(drawing, 1494, 1494, 4095, 4095, 0),
		(drawing, 1495, 1495, 4095, 4095, 0),
		(drawing, 1496, 1496, 4095, 4095, 0),
		(drawing, 1497, 1497, 4095, 4095, 0),
		(drawing, 1498, 1498, 4095, 4095, 0),
		(drawing, 1499, 1499, 4095, 4095, 0),
		(drawing, 1500, 1500, 4095, 4095, 0),
		(drawing, 1501, 1501, 4095, 4095, 0),
		(drawing, 1502, 1502, 4095, 4095, 0),
		(drawing, 1503, 1503, 4095, 4095, 0),
		(drawing, 1504, 1504, 4095, 4095, 0),
		(drawing, 1505, 1505, 4095, 4095, 0),
		(drawing, 1506, 1506, 4095, 4095, 0),
		(drawing, 1507, 1507, 4095, 4095, 0),
		(drawing, 1508, 1508, 4095, 4095, 0),
		(drawing, 1509, 1509, 4095, 4095, 0),
		(drawing, 1510, 1510, 4095, 4095, 0),
		(drawing, 1511, 1511, 4095, 4095, 0),
		(drawing, 1512, 1512, 4095, 4095, 0),
		(drawing, 1513, 1513, 4095, 4095, 0),
		(drawing, 1514, 1514, 4095, 4095, 0),
		(drawing, 1515, 1515, 4095, 4095, 0),
		(drawing, 1516, 1516, 4095, 4095, 0),
		(drawing, 1517, 1517, 4095, 4095, 0),
		(drawing, 1518, 1518, 4095, 4095, 0),
		(drawing, 1519, 1519, 4095, 4095, 0),
		(drawing, 1520, 1520, 4095, 4095, 0),
		(drawing, 1521, 1521, 4095, 4095, 0),
		(drawing, 1522, 1522, 4095, 4095, 0),
		(drawing, 1523, 1523, 4095, 4095, 0),
		(drawing, 1524, 1524, 4095, 4095, 0),
		(drawing, 1525, 1525, 4095, 4095, 0),
		(drawing, 1526, 1526, 4095, 4095, 0),
		(drawing, 1527, 1527, 4095, 4095, 0),
		(drawing, 1528, 1528, 4095, 4095, 0),
		(drawing, 1529, 1529, 4095, 4095, 0),
		(drawing, 1530, 1530, 4095, 4095, 0),
		(drawing, 1531, 1531, 4095, 4095, 0),
		(drawing, 1532, 1532, 4095, 4095, 0),
		(drawing, 1533, 1533, 4095, 4095, 0),
		(drawing, 1534, 1534, 4095, 4095, 0),
		(drawing, 1535, 1535, 4095, 4095, 0),
		(drawing, 1536, 1536, 4095, 4095, 0),
		(drawing, 1537, 1537, 4095, 4095, 0),
		(drawing, 1538, 1538, 4095, 4095, 0),
		(drawing, 1539, 1539, 4095, 4095, 0),
		(drawing, 1540, 1540, 4095, 4095, 0),
		(drawing, 1541, 1541, 4095, 4095, 0),
		(drawing, 1542, 1542, 4095, 4095, 0),
		(drawing, 1543, 1543, 4095, 4095, 0),
		(drawing, 1544, 1544, 4095, 4095, 0),
		(drawing, 1545, 1545, 4095, 4095, 0),
		(drawing, 1546, 1546, 4095, 4095, 0),
		(drawing, 1547, 1547, 4095, 4095, 0),
		(drawing, 1548, 1548, 4095, 4095, 0),
		(drawing, 1549, 1549, 4095, 4095, 0),
		(drawing, 1550, 1550, 4095, 4095, 0),
		(drawing, 1551, 1551, 4095, 4095, 0),
		(drawing, 1552, 1552, 4095, 4095, 0),
		(drawing, 1553, 1553, 4095, 4095, 0),
		(drawing, 1554, 1554, 4095, 4095, 0),
		(drawing, 1555, 1555, 4095, 4095, 0),
		(drawing, 1556, 1556, 4095, 4095, 0),
		(drawing, 1557, 1557, 4095, 4095, 0),
		(drawing, 1558, 1558, 4095, 4095, 0),
		(drawing, 1559, 1559, 4095, 4095, 0),
		(drawing, 1560, 1560, 4095, 4095, 0),
		(drawing, 1561, 1561, 4095, 4095, 0),
		(drawing, 1562, 1562, 4095, 4095, 0),
		(drawing, 1563, 1563, 4095, 4095, 0),
		(drawing, 1564, 1564, 4095, 4095, 0),
		(drawing, 1565, 1565, 4095, 4095, 0),
		(drawing, 1566, 1566, 4095, 4095, 0),
		(drawing, 1567, 1567, 4095, 4095, 0),
		(drawing, 1568, 1568, 4095, 4095, 0),
		(drawing, 1569, 1569, 4095, 4095, 0),
		(drawing, 1570, 1570, 4095, 4095, 0),
		(drawing, 1571, 1571, 4095, 4095, 0),
		(drawing, 1572, 1572, 4095, 4095, 0),
		(drawing, 1573, 1573, 4095, 4095, 0),
		(drawing, 1574, 1574, 4095, 4095, 0),
		(drawing, 1575, 1575, 4095, 4095, 0),
		(drawing, 1576, 1576, 4095, 4095, 0),
		(drawing, 1577, 1577, 4095, 4095, 0),
		(drawing, 1578, 1578, 4095, 4095, 0),
		(drawing, 1579, 1579, 4095, 4095, 0),
		(drawing, 1580, 1580, 4095, 4095, 0),
		(drawing, 1581, 1581, 4095, 4095, 0),
		(drawing, 1582, 1582, 4095, 4095, 0),
		(drawing, 1583, 1583, 4095, 4095, 0),
		(drawing, 1584, 1584, 4095, 4095, 0),
		(drawing, 1585, 1585, 4095, 4095, 0),
		(drawing, 1586, 1586, 4095, 4095, 0),
		(drawing, 1587, 1587, 4095, 4095, 0),
		(drawing, 1588, 1588, 4095, 4095, 0),
		(drawing, 1589, 1589, 4095, 4095, 0),
		(drawing, 1590, 1590, 4095, 4095, 0),
		(drawing, 1591, 1591, 4095, 4095, 0),
		(drawing, 1592, 1592, 4095, 4095, 0),
		(drawing, 1593, 1593, 4095, 4095, 0),
		(drawing, 1594, 1594, 4095, 4095, 0),
		(drawing, 1595, 1595, 4095, 4095, 0),
		(drawing, 1596, 1596, 4095, 4095, 0),
		(drawing, 1597, 1597, 4095, 4095, 0),
		(drawing, 1598, 1598, 4095, 4095, 0),
		(drawing, 1599, 1599, 4095, 4095, 0),
		(drawing, 1600, 1600, 4095, 4095, 0),
		(drawing, 1601, 1601, 4095, 4095, 0),
		(drawing, 1602, 1602, 4095, 4095, 0),
		(drawing, 1603, 1603, 4095, 4095, 0),
		(drawing, 1604, 1604, 4095, 4095, 0),
		(drawing, 1605, 1605, 4095, 4095, 0),
		(drawing, 1606, 1606, 4095, 4095, 0),
		(drawing, 1607, 1607, 4095, 4095, 0),
		(drawing, 1608, 1608, 4095, 4095, 0),
		(drawing, 1609, 1609, 4095, 4095, 0),
		(drawing, 1610, 1610, 4095, 4095, 0),
		(drawing, 1611, 1611, 4095, 4095, 0),
		(drawing, 1612, 1612, 4095, 4095, 0),
		(drawing, 1613, 1613, 4095, 4095, 0),
		(drawing, 1614, 1614, 4095, 4095, 0),
		(drawing, 1615, 1615, 4095, 4095, 0),
		(drawing, 1616, 1616, 4095, 4095, 0),
		(drawing, 1617, 1617, 4095, 4095, 0),
		(drawing, 1618, 1618, 4095, 4095, 0),
		(drawing, 1619, 1619, 4095, 4095, 0),
		(drawing, 1620, 1620, 4095, 4095, 0),
		(drawing, 1621, 1621, 4095, 4095, 0),
		(drawing, 1622, 1622, 4095, 4095, 0),
		(drawing, 1623, 1623, 4095, 4095, 0),
		(drawing, 1624, 1624, 4095, 4095, 0),
		(drawing, 1625, 1625, 4095, 4095, 0),
		(drawing, 1626, 1626, 4095, 4095, 0),
		(drawing, 1627, 1627, 4095, 4095, 0),
		(drawing, 1628, 1628, 4095, 4095, 0),
		(drawing, 1629, 1629, 4095, 4095, 0),
		(drawing, 1630, 1630, 4095, 4095, 0),
		(drawing, 1631, 1631, 4095, 4095, 0),
		(drawing, 1632, 1632, 4095, 4095, 0),
		(drawing, 1633, 1633, 4095, 4095, 0),
		(drawing, 1634, 1634, 4095, 4095, 0),
		(drawing, 1635, 1635, 4095, 4095, 0),
		(drawing, 1636, 1636, 4095, 4095, 0),
		(drawing, 1637, 1637, 4095, 4095, 0),
		(drawing, 1638, 1638, 4095, 4095, 0),
		(drawing, 1639, 1639, 4095, 4095, 0),
		(drawing, 1640, 1640, 4095, 4095, 0),
		(drawing, 1641, 1641, 4095, 4095, 0),
		(drawing, 1642, 1642, 4095, 4095, 0),
		(drawing, 1643, 1643, 4095, 4095, 0),
		(drawing, 1644, 1644, 4095, 4095, 0),
		(drawing, 1645, 1645, 4095, 4095, 0),
		(drawing, 1646, 1646, 4095, 4095, 0),
		(drawing, 1647, 1647, 4095, 4095, 0),
		(drawing, 1648, 1648, 4095, 4095, 0),
		(drawing, 1649, 1649, 4095, 4095, 0),
		(drawing, 1650, 1650, 4095, 4095, 0),
		(drawing, 1651, 1651, 4095, 4095, 0),
		(drawing, 1652, 1652, 4095, 4095, 0),
		(drawing, 1653, 1653, 4095, 4095, 0),
		(drawing, 1654, 1654, 4095, 4095, 0),
		(drawing, 1655, 1655, 4095, 4095, 0),
		(drawing, 1656, 1656, 4095, 4095, 0),
		(drawing, 1657, 1657, 4095, 4095, 0),
		(drawing, 1658, 1658, 4095, 4095, 0),
		(drawing, 1659, 1659, 4095, 4095, 0),
		(drawing, 1660, 1660, 4095, 4095, 0),
		(drawing, 1661, 1661, 4095, 4095, 0),
		(drawing, 1662, 1662, 4095, 4095, 0),
		(drawing, 1663, 1663, 4095, 4095, 0),
		(drawing, 1664, 1664, 4095, 4095, 0),
		(drawing, 1665, 1665, 4095, 4095, 0),
		(drawing, 1666, 1666, 4095, 4095, 0),
		(drawing, 1667, 1667, 4095, 4095, 0),
		(drawing, 1668, 1668, 4095, 4095, 0),
		(drawing, 1669, 1669, 4095, 4095, 0),
		(drawing, 1670, 1670, 4095, 4095, 0),
		(drawing, 1671, 1671, 4095, 4095, 0),
		(drawing, 1672, 1672, 4095, 4095, 0),
		(drawing, 1673, 1673, 4095, 4095, 0),
		(drawing, 1674, 1674, 4095, 4095, 0),
		(drawing, 1675, 1675, 4095, 4095, 0),
		(drawing, 1676, 1676, 4095, 4095, 0),
		(drawing, 1677, 1677, 4095, 4095, 0),
		(drawing, 1678, 1678, 4095, 4095, 0),
		(drawing, 1679, 1679, 4095, 4095, 0),
		(drawing, 1680, 1680, 4095, 4095, 0),
		(drawing, 1681, 1681, 4095, 4095, 0),
		(drawing, 1682, 1682, 4095, 4095, 0),
		(drawing, 1683, 1683, 4095, 4095, 0),
		(drawing, 1684, 1684, 4095, 4095, 0),
		(drawing, 1685, 1685, 4095, 4095, 0),
		(drawing, 1686, 1686, 4095, 4095, 0),
		(drawing, 1687, 1687, 4095, 4095, 0),
		(drawing, 1688, 1688, 4095, 4095, 0),
		(drawing, 1689, 1689, 4095, 4095, 0),
		(drawing, 1690, 1690, 4095, 4095, 0),
		(drawing, 1691, 1691, 4095, 4095, 0),
		(drawing, 1692, 1692, 4095, 4095, 0),
		(drawing, 1693, 1693, 4095, 4095, 0),
		(drawing, 1694, 1694, 4095, 4095, 0),
		(drawing, 1695, 1695, 4095, 4095, 0),
		(drawing, 1696, 1696, 4095, 4095, 0),
		(drawing, 1697, 1697, 4095, 4095, 0),
		(drawing, 1698, 1698, 4095, 4095, 0),
		(drawing, 1699, 1699, 4095, 4095, 0),
		(drawing, 1700, 1700, 4095, 4095, 0),
		(drawing, 1701, 1701, 4095, 4095, 0),
		(drawing, 1702, 1702, 4095, 4095, 0),
		(drawing, 1703, 1703, 4095, 4095, 0),
		(drawing, 1704, 1704, 4095, 4095, 0),
		(drawing, 1705, 1705, 4095, 4095, 0),
		(drawing, 1706, 1706, 4095, 4095, 0),
		(drawing, 1707, 1707, 4095, 4095, 0),
		(drawing, 1708, 1708, 4095, 4095, 0),
		(drawing, 1709, 1709, 4095, 4095, 0),
		(drawing, 1710, 1710, 4095, 4095, 0),
		(drawing, 1711, 1711, 4095, 4095, 0),
		(drawing, 1712, 1712, 4095, 4095, 0),
		(drawing, 1713, 1713, 4095, 4095, 0),
		(drawing, 1714, 1714, 4095, 4095, 0),
		(drawing, 1715, 1715, 4095, 4095, 0),
		(drawing, 1716, 1716, 4095, 4095, 0),
		(drawing, 1717, 1717, 4095, 4095, 0),
		(drawing, 1718, 1718, 4095, 4095, 0),
		(drawing, 1719, 1719, 4095, 4095, 0),
		(drawing, 1720, 1720, 4095, 4095, 0),
		(drawing, 1721, 1721, 4095, 4095, 0),
		(drawing, 1722, 1722, 4095, 4095, 0),
		(drawing, 1723, 1723, 4095, 4095, 0),
		(drawing, 1724, 1724, 4095, 4095, 0),
		(drawing, 1725, 1725, 4095, 4095, 0),
		(drawing, 1726, 1726, 4095, 4095, 0),
		(drawing, 1727, 1727, 4095, 4095, 0),
		(drawing, 1728, 1728, 4095, 4095, 0),
		(drawing, 1729, 1729, 4095, 4095, 0),
		(drawing, 1730, 1730, 4095, 4095, 0),
		(drawing, 1731, 1731, 4095, 4095, 0),
		(drawing, 1732, 1732, 4095, 4095, 0),
		(drawing, 1733, 1733, 4095, 4095, 0),
		(drawing, 1734, 1734, 4095, 4095, 0),
		(drawing, 1735, 1735, 4095, 4095, 0),
		(drawing, 1736, 1736, 4095, 4095, 0),
		(drawing, 1737, 1737, 4095, 4095, 0),
		(drawing, 1738, 1738, 4095, 4095, 0),
		(drawing, 1739, 1739, 4095, 4095, 0),
		(drawing, 1740, 1740, 4095, 4095, 0),
		(drawing, 1741, 1741, 4095, 4095, 0),
		(drawing, 1742, 1742, 4095, 4095, 0),
		(drawing, 1743, 1743, 4095, 4095, 0),
		(drawing, 1744, 1744, 4095, 4095, 0),
		(drawing, 1745, 1745, 4095, 4095, 0),
		(drawing, 1746, 1746, 4095, 4095, 0),
		(drawing, 1747, 1747, 4095, 4095, 0),
		(drawing, 1748, 1748, 4095, 4095, 0),
		(drawing, 1749, 1749, 4095, 4095, 0),
		(drawing, 1750, 1750, 4095, 4095, 0),
		(drawing, 1751, 1751, 4095, 4095, 0),
		(drawing, 1752, 1752, 4095, 4095, 0),
		(drawing, 1753, 1753, 4095, 4095, 0),
		(drawing, 1754, 1754, 4095, 4095, 0),
		(drawing, 1755, 1755, 4095, 4095, 0),
		(drawing, 1756, 1756, 4095, 4095, 0),
		(drawing, 1757, 1757, 4095, 4095, 0),
		(drawing, 1758, 1758, 4095, 4095, 0),
		(drawing, 1759, 1759, 4095, 4095, 0),
		(drawing, 1760, 1760, 4095, 4095, 0),
		(drawing, 1761, 1761, 4095, 4095, 0),
		(drawing, 1762, 1762, 4095, 4095, 0),
		(drawing, 1763, 1763, 4095, 4095, 0),
		(drawing, 1764, 1764, 4095, 4095, 0),
		(drawing, 1765, 1765, 4095, 4095, 0),
		(drawing, 1766, 1766, 4095, 4095, 0),
		(drawing, 1767, 1767, 4095, 4095, 0),
		(drawing, 1768, 1768, 4095, 4095, 0),
		(drawing, 1769, 1769, 4095, 4095, 0),
		(drawing, 1770, 1770, 4095, 4095, 0),
		(drawing, 1771, 1771, 4095, 4095, 0),
		(drawing, 1772, 1772, 4095, 4095, 0),
		(drawing, 1773, 1773, 4095, 4095, 0),
		(drawing, 1774, 1774, 4095, 4095, 0),
		(drawing, 1775, 1775, 4095, 4095, 0),
		(drawing, 1776, 1776, 4095, 4095, 0),
		(drawing, 1777, 1777, 4095, 4095, 0),
		(drawing, 1778, 1778, 4095, 4095, 0),
		(drawing, 1779, 1779, 4095, 4095, 0),
		(drawing, 1780, 1780, 4095, 4095, 0),
		(drawing, 1781, 1781, 4095, 4095, 0),
		(drawing, 1782, 1782, 4095, 4095, 0),
		(drawing, 1783, 1783, 4095, 4095, 0),
		(drawing, 1784, 1784, 4095, 4095, 0),
		(drawing, 1785, 1785, 4095, 4095, 0),
		(drawing, 1786, 1786, 4095, 4095, 0),
		(drawing, 1787, 1787, 4095, 4095, 0),
		(drawing, 1788, 1788, 4095, 4095, 0),
		(drawing, 1789, 1789, 4095, 4095, 0),
		(drawing, 1790, 1790, 4095, 4095, 0),
		(drawing, 1791, 1791, 4095, 4095, 0),
		(drawing, 1792, 1792, 4095, 4095, 0),
		(drawing, 1793, 1793, 4095, 4095, 0),
		(drawing, 1794, 1794, 4095, 4095, 0),
		(drawing, 1795, 1795, 4095, 4095, 0),
		(drawing, 1796, 1796, 4095, 4095, 0),
		(drawing, 1797, 1797, 4095, 4095, 0),
		(drawing, 1798, 1798, 4095, 4095, 0),
		(drawing, 1799, 1799, 4095, 4095, 0),
		(drawing, 1800, 1800, 4095, 4095, 0),
		(drawing, 1801, 1801, 4095, 4095, 0),
		(drawing, 1802, 1802, 4095, 4095, 0),
		(drawing, 1803, 1803, 4095, 4095, 0),
		(drawing, 1804, 1804, 4095, 4095, 0),
		(drawing, 1805, 1805, 4095, 4095, 0),
		(drawing, 1806, 1806, 4095, 4095, 0),
		(drawing, 1807, 1807, 4095, 4095, 0),
		(drawing, 1808, 1808, 4095, 4095, 0),
		(drawing, 1809, 1809, 4095, 4095, 0),
		(drawing, 1810, 1810, 4095, 4095, 0),
		(drawing, 1811, 1811, 4095, 4095, 0),
		(drawing, 1812, 1812, 4095, 4095, 0),
		(drawing, 1813, 1813, 4095, 4095, 0),
		(drawing, 1814, 1814, 4095, 4095, 0),
		(drawing, 1815, 1815, 4095, 4095, 0),
		(drawing, 1816, 1816, 4095, 4095, 0),
		(drawing, 1817, 1817, 4095, 4095, 0),
		(drawing, 1818, 1818, 4095, 4095, 0),
		(drawing, 1819, 1819, 4095, 4095, 0),
		(drawing, 1820, 1820, 4095, 4095, 0),
		(drawing, 1821, 1821, 4095, 4095, 0),
		(drawing, 1822, 1822, 4095, 4095, 0),
		(drawing, 1823, 1823, 4095, 4095, 0),
		(drawing, 1824, 1824, 4095, 4095, 0),
		(drawing, 1825, 1825, 4095, 4095, 0),
		(drawing, 1826, 1826, 4095, 4095, 0),
		(drawing, 1827, 1827, 4095, 4095, 0),
		(drawing, 1828, 1828, 4095, 4095, 0),
		(drawing, 1829, 1829, 4095, 4095, 0),
		(drawing, 1830, 1830, 4095, 4095, 0),
		(drawing, 1831, 1831, 4095, 4095, 0),
		(drawing, 1832, 1832, 4095, 4095, 0),
		(drawing, 1833, 1833, 4095, 4095, 0),
		(drawing, 1834, 1834, 4095, 4095, 0),
		(drawing, 1835, 1835, 4095, 4095, 0),
		(drawing, 1836, 1836, 4095, 4095, 0),
		(drawing, 1837, 1837, 4095, 4095, 0),
		(drawing, 1838, 1838, 4095, 4095, 0),
		(drawing, 1839, 1839, 4095, 4095, 0),
		(drawing, 1840, 1840, 4095, 4095, 0),
		(drawing, 1841, 1841, 4095, 4095, 0),
		(drawing, 1842, 1842, 4095, 4095, 0),
		(drawing, 1843, 1843, 4095, 4095, 0),
		(drawing, 1844, 1844, 4095, 4095, 0),
		(drawing, 1845, 1845, 4095, 4095, 0),
		(drawing, 1846, 1846, 4095, 4095, 0),
		(drawing, 1847, 1847, 4095, 4095, 0),
		(drawing, 1848, 1848, 4095, 4095, 0),
		(drawing, 1849, 1849, 4095, 4095, 0),
		(drawing, 1850, 1850, 4095, 4095, 0),
		(drawing, 1851, 1851, 4095, 4095, 0),
		(drawing, 1852, 1852, 4095, 4095, 0),
		(drawing, 1853, 1853, 4095, 4095, 0),
		(drawing, 1854, 1854, 4095, 4095, 0),
		(drawing, 1855, 1855, 4095, 4095, 0),
		(drawing, 1856, 1856, 4095, 4095, 0),
		(drawing, 1857, 1857, 4095, 4095, 0),
		(drawing, 1858, 1858, 4095, 4095, 0),
		(drawing, 1859, 1859, 4095, 4095, 0),
		(drawing, 1860, 1860, 4095, 4095, 0),
		(drawing, 1861, 1861, 4095, 4095, 0),
		(drawing, 1862, 1862, 4095, 4095, 0),
		(drawing, 1863, 1863, 4095, 4095, 0),
		(drawing, 1864, 1864, 4095, 4095, 0),
		(drawing, 1865, 1865, 4095, 4095, 0),
		(drawing, 1866, 1866, 4095, 4095, 0),
		(drawing, 1867, 1867, 4095, 4095, 0),
		(drawing, 1868, 1868, 4095, 4095, 0),
		(drawing, 1869, 1869, 4095, 4095, 0),
		(drawing, 1870, 1870, 4095, 4095, 0),
		(drawing, 1871, 1871, 4095, 4095, 0),
		(drawing, 1872, 1872, 4095, 4095, 0),
		(drawing, 1873, 1873, 4095, 4095, 0),
		(drawing, 1874, 1874, 4095, 4095, 0),
		(drawing, 1875, 1875, 4095, 4095, 0),
		(drawing, 1876, 1876, 4095, 4095, 0),
		(drawing, 1877, 1877, 4095, 4095, 0),
		(drawing, 1878, 1878, 4095, 4095, 0),
		(drawing, 1879, 1879, 4095, 4095, 0),
		(drawing, 1880, 1880, 4095, 4095, 0),
		(drawing, 1881, 1881, 4095, 4095, 0),
		(drawing, 1882, 1882, 4095, 4095, 0),
		(drawing, 1883, 1883, 4095, 4095, 0),
		(drawing, 1884, 1884, 4095, 4095, 0),
		(drawing, 1885, 1885, 4095, 4095, 0),
		(drawing, 1886, 1886, 4095, 4095, 0),
		(drawing, 1887, 1887, 4095, 4095, 0),
		(drawing, 1888, 1888, 4095, 4095, 0),
		(drawing, 1889, 1889, 4095, 4095, 0),
		(drawing, 1890, 1890, 4095, 4095, 0),
		(drawing, 1891, 1891, 4095, 4095, 0),
		(drawing, 1892, 1892, 4095, 4095, 0),
		(drawing, 1893, 1893, 4095, 4095, 0),
		(drawing, 1894, 1894, 4095, 4095, 0),
		(drawing, 1895, 1895, 4095, 4095, 0),
		(drawing, 1896, 1896, 4095, 4095, 0),
		(drawing, 1897, 1897, 4095, 4095, 0),
		(drawing, 1898, 1898, 4095, 4095, 0),
		(drawing, 1899, 1899, 4095, 4095, 0),
		(drawing, 1900, 1900, 4095, 4095, 0),
		(drawing, 1901, 1901, 4095, 4095, 0),
		(drawing, 1902, 1902, 4095, 4095, 0),
		(drawing, 1903, 1903, 4095, 4095, 0),
		(drawing, 1904, 1904, 4095, 4095, 0),
		(drawing, 1905, 1905, 4095, 4095, 0),
		(drawing, 1906, 1906, 4095, 4095, 0),
		(drawing, 1907, 1907, 4095, 4095, 0),
		(drawing, 1908, 1908, 4095, 4095, 0),
		(drawing, 1909, 1909, 4095, 4095, 0),
		(drawing, 1910, 1910, 4095, 4095, 0),
		(drawing, 1911, 1911, 4095, 4095, 0),
		(drawing, 1912, 1912, 4095, 4095, 0),
		(drawing, 1913, 1913, 4095, 4095, 0),
		(drawing, 1914, 1914, 4095, 4095, 0),
		(drawing, 1915, 1915, 4095, 4095, 0),
		(drawing, 1916, 1916, 4095, 4095, 0),
		(drawing, 1917, 1917, 4095, 4095, 0),
		(drawing, 1918, 1918, 4095, 4095, 0),
		(drawing, 1919, 1919, 4095, 4095, 0),
		(drawing, 1920, 1920, 4095, 4095, 0),
		(drawing, 1921, 1921, 4095, 4095, 0),
		(drawing, 1922, 1922, 4095, 4095, 0),
		(drawing, 1923, 1923, 4095, 4095, 0),
		(drawing, 1924, 1924, 4095, 4095, 0),
		(drawing, 1925, 1925, 4095, 4095, 0),
		(drawing, 1926, 1926, 4095, 4095, 0),
		(drawing, 1927, 1927, 4095, 4095, 0),
		(drawing, 1928, 1928, 4095, 4095, 0),
		(drawing, 1929, 1929, 4095, 4095, 0),
		(drawing, 1930, 1930, 4095, 4095, 0),
		(drawing, 1931, 1931, 4095, 4095, 0),
		(drawing, 1932, 1932, 4095, 4095, 0),
		(drawing, 1933, 1933, 4095, 4095, 0),
		(drawing, 1934, 1934, 4095, 4095, 0),
		(drawing, 1935, 1935, 4095, 4095, 0),
		(drawing, 1936, 1936, 4095, 4095, 0),
		(drawing, 1937, 1937, 4095, 4095, 0),
		(drawing, 1938, 1938, 4095, 4095, 0),
		(drawing, 1939, 1939, 4095, 4095, 0),
		(drawing, 1940, 1940, 4095, 4095, 0),
		(drawing, 1941, 1941, 4095, 4095, 0),
		(drawing, 1942, 1942, 4095, 4095, 0),
		(drawing, 1943, 1943, 4095, 4095, 0),
		(drawing, 1944, 1944, 4095, 4095, 0),
		(drawing, 1945, 1945, 4095, 4095, 0),
		(drawing, 1946, 1946, 4095, 4095, 0),
		(drawing, 1947, 1947, 4095, 4095, 0),
		(drawing, 1948, 1948, 4095, 4095, 0),
		(drawing, 1949, 1949, 4095, 4095, 0),
		(drawing, 1950, 1950, 4095, 4095, 0),
		(drawing, 1951, 1951, 4095, 4095, 0),
		(drawing, 1952, 1952, 4095, 4095, 0),
		(drawing, 1953, 1953, 4095, 4095, 0),
		(drawing, 1954, 1954, 4095, 4095, 0),
		(drawing, 1955, 1955, 4095, 4095, 0),
		(drawing, 1956, 1956, 4095, 4095, 0),
		(drawing, 1957, 1957, 4095, 4095, 0),
		(drawing, 1958, 1958, 4095, 4095, 0),
		(drawing, 1959, 1959, 4095, 4095, 0),
		(drawing, 1960, 1960, 4095, 4095, 0),
		(drawing, 1961, 1961, 4095, 4095, 0),
		(drawing, 1962, 1962, 4095, 4095, 0),
		(drawing, 1963, 1963, 4095, 4095, 0),
		(drawing, 1964, 1964, 4095, 4095, 0),
		(drawing, 1965, 1965, 4095, 4095, 0),
		(drawing, 1966, 1966, 4095, 4095, 0),
		(drawing, 1967, 1967, 4095, 4095, 0),
		(drawing, 1968, 1968, 4095, 4095, 0),
		(drawing, 1969, 1969, 4095, 4095, 0),
		(drawing, 1970, 1970, 4095, 4095, 0),
		(drawing, 1971, 1971, 4095, 4095, 0),
		(drawing, 1972, 1972, 4095, 4095, 0),
		(drawing, 1973, 1973, 4095, 4095, 0),
		(drawing, 1974, 1974, 4095, 4095, 0),
		(drawing, 1975, 1975, 4095, 4095, 0),
		(drawing, 1976, 1976, 4095, 4095, 0),
		(drawing, 1977, 1977, 4095, 4095, 0),
		(drawing, 1978, 1978, 4095, 4095, 0),
		(drawing, 1979, 1979, 4095, 4095, 0),
		(drawing, 1980, 1980, 4095, 4095, 0),
		(drawing, 1981, 1981, 4095, 4095, 0),
		(drawing, 1982, 1982, 4095, 4095, 0),
		(drawing, 1983, 1983, 4095, 4095, 0),
		(drawing, 1984, 1984, 4095, 4095, 0),
		(drawing, 1985, 1985, 4095, 4095, 0),
		(drawing, 1986, 1986, 4095, 4095, 0),
		(drawing, 1987, 1987, 4095, 4095, 0),
		(drawing, 1988, 1988, 4095, 4095, 0),
		(drawing, 1989, 1989, 4095, 4095, 0),
		(drawing, 1990, 1990, 4095, 4095, 0),
		(drawing, 1991, 1991, 4095, 4095, 0),
		(drawing, 1992, 1992, 4095, 4095, 0),
		(drawing, 1993, 1993, 4095, 4095, 0),
		(drawing, 1994, 1994, 4095, 4095, 0),
		(drawing, 1995, 1995, 4095, 4095, 0),
		(drawing, 1996, 1996, 4095, 4095, 0),
		(drawing, 1997, 1997, 4095, 4095, 0),
		(drawing, 1998, 1998, 4095, 4095, 0),
		(drawing, 1999, 1999, 4095, 4095, 0),
		(drawing, 2000, 2000, 4095, 4095, 0),
		(drawing, 2001, 2001, 4095, 4095, 0),
		(drawing, 2002, 2002, 4095, 4095, 0),
		(drawing, 2003, 2003, 4095, 4095, 0),
		(drawing, 2004, 2004, 4095, 4095, 0),
		(drawing, 2005, 2005, 4095, 4095, 0),
		(drawing, 2006, 2006, 4095, 4095, 0),
		(drawing, 2007, 2007, 4095, 4095, 0),
		(drawing, 2008, 2008, 4095, 4095, 0),
		(drawing, 2009, 2009, 4095, 4095, 0),
		(drawing, 2010, 2010, 4095, 4095, 0),
		(drawing, 2011, 2011, 4095, 4095, 0),
		(drawing, 2012, 2012, 4095, 4095, 0),
		(drawing, 2013, 2013, 4095, 4095, 0),
		(drawing, 2014, 2014, 4095, 4095, 0),
		(drawing, 2015, 2015, 4095, 4095, 0),
		(drawing, 2016, 2016, 4095, 4095, 0),
		(drawing, 2017, 2017, 4095, 4095, 0),
		(drawing, 2018, 2018, 4095, 4095, 0),
		(drawing, 2019, 2019, 4095, 4095, 0),
		(drawing, 2020, 2020, 4095, 4095, 0),
		(drawing, 2021, 2021, 4095, 4095, 0),
		(drawing, 2022, 2022, 4095, 4095, 0),
		(drawing, 2023, 2023, 4095, 4095, 0),
		(drawing, 2024, 2024, 4095, 4095, 0),
		(drawing, 2025, 2025, 4095, 4095, 0),
		(drawing, 2026, 2026, 4095, 4095, 0),
		(drawing, 2027, 2027, 4095, 4095, 0),
		(drawing, 2028, 2028, 4095, 4095, 0),
		(drawing, 2029, 2029, 4095, 4095, 0),
		(drawing, 2030, 2030, 4095, 4095, 0),
		(drawing, 2031, 2031, 4095, 4095, 0),
		(drawing, 2032, 2032, 4095, 4095, 0),
		(drawing, 2033, 2033, 4095, 4095, 0),
		(drawing, 2034, 2034, 4095, 4095, 0),
		(drawing, 2035, 2035, 4095, 4095, 0),
		(drawing, 2036, 2036, 4095, 4095, 0),
		(drawing, 2037, 2037, 4095, 4095, 0),
		(drawing, 2038, 2038, 4095, 4095, 0),
		(drawing, 2039, 2039, 4095, 4095, 0),
		(drawing, 2040, 2040, 4095, 4095, 0),
		(drawing, 2041, 2041, 4095, 4095, 0),
		(drawing, 2042, 2042, 4095, 4095, 0),
		(drawing, 2043, 2043, 4095, 4095, 0),
		(drawing, 2044, 2044, 4095, 4095, 0),
		(drawing, 2045, 2045, 4095, 4095, 0),
		(drawing, 2046, 2046, 4095, 4095, 0),
		(drawing, 2047, 2047, 4095, 4095, 0),
		(drawing, 2048, 2048, 4095, 4095, 0),
		(drawing, 2049, 2049, 4095, 4095, 0),
		(drawing, 2050, 2050, 4095, 4095, 0),
		(drawing, 2051, 2051, 4095, 4095, 0),
		(drawing, 2052, 2052, 4095, 4095, 0),
		(drawing, 2053, 2053, 4095, 4095, 0),
		(drawing, 2054, 2054, 4095, 4095, 0),
		(drawing, 2055, 2055, 4095, 4095, 0),
		(drawing, 2056, 2056, 4095, 4095, 0),
		(drawing, 2057, 2057, 4095, 4095, 0),
		(drawing, 2058, 2058, 4095, 4095, 0),
		(drawing, 2059, 2059, 4095, 4095, 0),
		(drawing, 2060, 2060, 4095, 4095, 0),
		(drawing, 2061, 2061, 4095, 4095, 0),
		(drawing, 2062, 2062, 4095, 4095, 0),
		(drawing, 2063, 2063, 4095, 4095, 0),
		(drawing, 2064, 2064, 4095, 4095, 0),
		(drawing, 2065, 2065, 4095, 4095, 0),
		(drawing, 2066, 2066, 4095, 4095, 0),
		(drawing, 2067, 2067, 4095, 4095, 0),
		(drawing, 2068, 2068, 4095, 4095, 0),
		(drawing, 2069, 2069, 4095, 4095, 0),
		(drawing, 2070, 2070, 4095, 4095, 0),
		(drawing, 2071, 2071, 4095, 4095, 0),
		(drawing, 2072, 2072, 4095, 4095, 0),
		(drawing, 2073, 2073, 4095, 4095, 0),
		(drawing, 2074, 2074, 4095, 4095, 0),
		(drawing, 2075, 2075, 4095, 4095, 0),
		(drawing, 2076, 2076, 4095, 4095, 0),
		(drawing, 2077, 2077, 4095, 4095, 0),
		(drawing, 2078, 2078, 4095, 4095, 0),
		(drawing, 2079, 2079, 4095, 4095, 0),
		(drawing, 2080, 2080, 4095, 4095, 0),
		(drawing, 2081, 2081, 4095, 4095, 0),
		(drawing, 2082, 2082, 4095, 4095, 0),
		(drawing, 2083, 2083, 4095, 4095, 0),
		(drawing, 2084, 2084, 4095, 4095, 0),
		(drawing, 2085, 2085, 4095, 4095, 0),
		(drawing, 2086, 2086, 4095, 4095, 0),
		(drawing, 2087, 2087, 4095, 4095, 0),
		(drawing, 2088, 2088, 4095, 4095, 0),
		(drawing, 2089, 2089, 4095, 4095, 0),
		(drawing, 2090, 2090, 4095, 4095, 0),
		(drawing, 2091, 2091, 4095, 4095, 0),
		(drawing, 2092, 2092, 4095, 4095, 0),
		(drawing, 2093, 2093, 4095, 4095, 0),
		(drawing, 2094, 2094, 4095, 4095, 0),
		(drawing, 2095, 2095, 4095, 4095, 0),
		(drawing, 2096, 2096, 4095, 4095, 0),
		(drawing, 2097, 2097, 4095, 4095, 0),
		(drawing, 2098, 2098, 4095, 4095, 0),
		(drawing, 2099, 2099, 4095, 4095, 0),
		(drawing, 2100, 2100, 4095, 4095, 0),
		(drawing, 2101, 2101, 4095, 4095, 0),
		(drawing, 2102, 2102, 4095, 4095, 0),
		(drawing, 2103, 2103, 4095, 4095, 0),
		(drawing, 2104, 2104, 4095, 4095, 0),
		(drawing, 2105, 2105, 4095, 4095, 0),
		(drawing, 2106, 2106, 4095, 4095, 0),
		(drawing, 2107, 2107, 4095, 4095, 0),
		(drawing, 2108, 2108, 4095, 4095, 0),
		(drawing, 2109, 2109, 4095, 4095, 0),
		(drawing, 2110, 2110, 4095, 4095, 0),
		(drawing, 2111, 2111, 4095, 4095, 0),
		(drawing, 2112, 2112, 4095, 4095, 0),
		(drawing, 2113, 2113, 4095, 4095, 0),
		(drawing, 2114, 2114, 4095, 4095, 0),
		(drawing, 2115, 2115, 4095, 4095, 0),
		(drawing, 2116, 2116, 4095, 4095, 0),
		(drawing, 2117, 2117, 4095, 4095, 0),
		(drawing, 2118, 2118, 4095, 4095, 0),
		(drawing, 2119, 2119, 4095, 4095, 0),
		(drawing, 2120, 2120, 4095, 4095, 0),
		(drawing, 2121, 2121, 4095, 4095, 0),
		(drawing, 2122, 2122, 4095, 4095, 0),
		(drawing, 2123, 2123, 4095, 4095, 0),
		(drawing, 2124, 2124, 4095, 4095, 0),
		(drawing, 2125, 2125, 4095, 4095, 0),
		(drawing, 2126, 2126, 4095, 4095, 0),
		(drawing, 2127, 2127, 4095, 4095, 0),
		(drawing, 2128, 2128, 4095, 4095, 0),
		(drawing, 2129, 2129, 4095, 4095, 0),
		(drawing, 2130, 2130, 4095, 4095, 0),
		(drawing, 2131, 2131, 4095, 4095, 0),
		(drawing, 2132, 2132, 4095, 4095, 0),
		(drawing, 2133, 2133, 4095, 4095, 0),
		(drawing, 2134, 2134, 4095, 4095, 0),
		(drawing, 2135, 2135, 4095, 4095, 0),
		(drawing, 2136, 2136, 4095, 4095, 0),
		(drawing, 2137, 2137, 4095, 4095, 0),
		(drawing, 2138, 2138, 4095, 4095, 0),
		(drawing, 2139, 2139, 4095, 4095, 0),
		(drawing, 2140, 2140, 4095, 4095, 0),
		(drawing, 2141, 2141, 4095, 4095, 0),
		(drawing, 2142, 2142, 4095, 4095, 0),
		(drawing, 2143, 2143, 4095, 4095, 0),
		(drawing, 2144, 2144, 4095, 4095, 0),
		(drawing, 2145, 2145, 4095, 4095, 0),
		(drawing, 2146, 2146, 4095, 4095, 0),
		(drawing, 2147, 2147, 4095, 4095, 0),
		(drawing, 2148, 2148, 4095, 4095, 0),
		(drawing, 2149, 2149, 4095, 4095, 0),
		(drawing, 2150, 2150, 4095, 4095, 0),
		(drawing, 2151, 2151, 4095, 4095, 0),
		(drawing, 2152, 2152, 4095, 4095, 0),
		(drawing, 2153, 2153, 4095, 4095, 0),
		(drawing, 2154, 2154, 4095, 4095, 0),
		(drawing, 2155, 2155, 4095, 4095, 0),
		(drawing, 2156, 2156, 4095, 4095, 0),
		(drawing, 2157, 2157, 4095, 4095, 0),
		(drawing, 2158, 2158, 4095, 4095, 0),
		(drawing, 2159, 2159, 4095, 4095, 0),
		(drawing, 2160, 2160, 4095, 4095, 0),
		(drawing, 2161, 2161, 4095, 4095, 0),
		(drawing, 2162, 2162, 4095, 4095, 0),
		(drawing, 2163, 2163, 4095, 4095, 0),
		(drawing, 2164, 2164, 4095, 4095, 0),
		(drawing, 2165, 2165, 4095, 4095, 0),
		(drawing, 2166, 2166, 4095, 4095, 0),
		(drawing, 2167, 2167, 4095, 4095, 0),
		(drawing, 2168, 2168, 4095, 4095, 0),
		(drawing, 2169, 2169, 4095, 4095, 0),
		(drawing, 2170, 2170, 4095, 4095, 0),
		(drawing, 2171, 2171, 4095, 4095, 0),
		(drawing, 2172, 2172, 4095, 4095, 0),
		(drawing, 2173, 2173, 4095, 4095, 0),
		(drawing, 2174, 2174, 4095, 4095, 0),
		(drawing, 2175, 2175, 4095, 4095, 0),
		(drawing, 2176, 2176, 4095, 4095, 0),
		(drawing, 2177, 2177, 4095, 4095, 0),
		(drawing, 2178, 2178, 4095, 4095, 0),
		(drawing, 2179, 2179, 4095, 4095, 0),
		(drawing, 2180, 2180, 4095, 4095, 0),
		(drawing, 2181, 2181, 4095, 4095, 0),
		(drawing, 2182, 2182, 4095, 4095, 0),
		(drawing, 2183, 2183, 4095, 4095, 0),
		(drawing, 2184, 2184, 4095, 4095, 0),
		(drawing, 2185, 2185, 4095, 4095, 0),
		(drawing, 2186, 2186, 4095, 4095, 0),
		(drawing, 2187, 2187, 4095, 4095, 0),
		(drawing, 2188, 2188, 4095, 4095, 0),
		(drawing, 2189, 2189, 4095, 4095, 0),
		(drawing, 2190, 2190, 4095, 4095, 0),
		(drawing, 2191, 2191, 4095, 4095, 0),
		(drawing, 2192, 2192, 4095, 4095, 0),
		(drawing, 2193, 2193, 4095, 4095, 0),
		(drawing, 2194, 2194, 4095, 4095, 0),
		(drawing, 2195, 2195, 4095, 4095, 0),
		(drawing, 2196, 2196, 4095, 4095, 0),
		(drawing, 2197, 2197, 4095, 4095, 0),
		(drawing, 2198, 2198, 4095, 4095, 0),
		(drawing, 2199, 2199, 4095, 4095, 0),
		(drawing, 2200, 2200, 4095, 4095, 0),
		(drawing, 2201, 2201, 4095, 4095, 0),
		(drawing, 2202, 2202, 4095, 4095, 0),
		(drawing, 2203, 2203, 4095, 4095, 0),
		(drawing, 2204, 2204, 4095, 4095, 0),
		(drawing, 2205, 2205, 4095, 4095, 0),
		(drawing, 2206, 2206, 4095, 4095, 0),
		(drawing, 2207, 2207, 4095, 4095, 0),
		(drawing, 2208, 2208, 4095, 4095, 0),
		(drawing, 2209, 2209, 4095, 4095, 0),
		(drawing, 2210, 2210, 4095, 4095, 0),
		(drawing, 2211, 2211, 4095, 4095, 0),
		(drawing, 2212, 2212, 4095, 4095, 0),
		(drawing, 2213, 2213, 4095, 4095, 0),
		(drawing, 2214, 2214, 4095, 4095, 0),
		(drawing, 2215, 2215, 4095, 4095, 0),
		(drawing, 2216, 2216, 4095, 4095, 0),
		(drawing, 2217, 2217, 4095, 4095, 0),
		(drawing, 2218, 2218, 4095, 4095, 0),
		(drawing, 2219, 2219, 4095, 4095, 0),
		(drawing, 2220, 2220, 4095, 4095, 0),
		(drawing, 2221, 2221, 4095, 4095, 0),
		(drawing, 2222, 2222, 4095, 4095, 0),
		(drawing, 2223, 2223, 4095, 4095, 0),
		(drawing, 2224, 2224, 4095, 4095, 0),
		(drawing, 2225, 2225, 4095, 4095, 0),
		(drawing, 2226, 2226, 4095, 4095, 0),
		(drawing, 2227, 2227, 4095, 4095, 0),
		(drawing, 2228, 2228, 4095, 4095, 0),
		(drawing, 2229, 2229, 4095, 4095, 0),
		(drawing, 2230, 2230, 4095, 4095, 0),
		(drawing, 2231, 2231, 4095, 4095, 0),
		(drawing, 2232, 2232, 4095, 4095, 0),
		(drawing, 2233, 2233, 4095, 4095, 0),
		(drawing, 2234, 2234, 4095, 4095, 0),
		(drawing, 2235, 2235, 4095, 4095, 0),
		(drawing, 2236, 2236, 4095, 4095, 0),
		(drawing, 2237, 2237, 4095, 4095, 0),
		(drawing, 2238, 2238, 4095, 4095, 0),
		(drawing, 2239, 2239, 4095, 4095, 0),
		(drawing, 2240, 2240, 4095, 4095, 0),
		(drawing, 2241, 2241, 4095, 4095, 0),
		(drawing, 2242, 2242, 4095, 4095, 0),
		(drawing, 2243, 2243, 4095, 4095, 0),
		(drawing, 2244, 2244, 4095, 4095, 0),
		(drawing, 2245, 2245, 4095, 4095, 0),
		(drawing, 2246, 2246, 4095, 4095, 0),
		(drawing, 2247, 2247, 4095, 4095, 0),
		(drawing, 2248, 2248, 4095, 4095, 0),
		(drawing, 2249, 2249, 4095, 4095, 0),
		(drawing, 2250, 2250, 4095, 4095, 0),
		(drawing, 2251, 2251, 4095, 4095, 0),
		(drawing, 2252, 2252, 4095, 4095, 0),
		(drawing, 2253, 2253, 4095, 4095, 0),
		(drawing, 2254, 2254, 4095, 4095, 0),
		(drawing, 2255, 2255, 4095, 4095, 0),
		(drawing, 2256, 2256, 4095, 4095, 0),
		(drawing, 2257, 2257, 4095, 4095, 0),
		(drawing, 2258, 2258, 4095, 4095, 0),
		(drawing, 2259, 2259, 4095, 4095, 0),
		(drawing, 2260, 2260, 4095, 4095, 0),
		(drawing, 2261, 2261, 4095, 4095, 0),
		(drawing, 2262, 2262, 4095, 4095, 0),
		(drawing, 2263, 2263, 4095, 4095, 0),
		(drawing, 2264, 2264, 4095, 4095, 0),
		(drawing, 2265, 2265, 4095, 4095, 0),
		(drawing, 2266, 2266, 4095, 4095, 0),
		(drawing, 2267, 2267, 4095, 4095, 0),
		(drawing, 2268, 2268, 4095, 4095, 0),
		(drawing, 2269, 2269, 4095, 4095, 0),
		(drawing, 2270, 2270, 4095, 4095, 0),
		(drawing, 2271, 2271, 4095, 4095, 0),
		(drawing, 2272, 2272, 4095, 4095, 0),
		(drawing, 2273, 2273, 4095, 4095, 0),
		(drawing, 2274, 2274, 4095, 4095, 0),
		(drawing, 2275, 2275, 4095, 4095, 0),
		(drawing, 2276, 2276, 4095, 4095, 0),
		(drawing, 2277, 2277, 4095, 4095, 0),
		(drawing, 2278, 2278, 4095, 4095, 0),
		(drawing, 2279, 2279, 4095, 4095, 0),
		(drawing, 2280, 2280, 4095, 4095, 0),
		(drawing, 2281, 2281, 4095, 4095, 0),
		(drawing, 2282, 2282, 4095, 4095, 0),
		(drawing, 2283, 2283, 4095, 4095, 0),
		(drawing, 2284, 2284, 4095, 4095, 0),
		(drawing, 2285, 2285, 4095, 4095, 0),
		(drawing, 2286, 2286, 4095, 4095, 0),
		(drawing, 2287, 2287, 4095, 4095, 0),
		(drawing, 2288, 2288, 4095, 4095, 0),
		(drawing, 2289, 2289, 4095, 4095, 0),
		(drawing, 2290, 2290, 4095, 4095, 0),
		(drawing, 2291, 2291, 4095, 4095, 0),
		(drawing, 2292, 2292, 4095, 4095, 0),
		(drawing, 2293, 2293, 4095, 4095, 0),
		(drawing, 2294, 2294, 4095, 4095, 0),
		(drawing, 2295, 2295, 4095, 4095, 0),
		(drawing, 2296, 2296, 4095, 4095, 0),
		(drawing, 2297, 2297, 4095, 4095, 0),
		(drawing, 2298, 2298, 4095, 4095, 0),
		(drawing, 2299, 2299, 4095, 4095, 0),
		(drawing, 2300, 2300, 4095, 4095, 0),
		(drawing, 2301, 2301, 4095, 4095, 0),
		(drawing, 2302, 2302, 4095, 4095, 0),
		(drawing, 2303, 2303, 4095, 4095, 0),
		(drawing, 2304, 2304, 4095, 4095, 0),
		(drawing, 2305, 2305, 4095, 4095, 0),
		(drawing, 2306, 2306, 4095, 4095, 0),
		(drawing, 2307, 2307, 4095, 4095, 0),
		(drawing, 2308, 2308, 4095, 4095, 0),
		(drawing, 2309, 2309, 4095, 4095, 0),
		(drawing, 2310, 2310, 4095, 4095, 0),
		(drawing, 2311, 2311, 4095, 4095, 0),
		(drawing, 2312, 2312, 4095, 4095, 0),
		(drawing, 2313, 2313, 4095, 4095, 0),
		(drawing, 2314, 2314, 4095, 4095, 0),
		(drawing, 2315, 2315, 4095, 4095, 0),
		(drawing, 2316, 2316, 4095, 4095, 0),
		(drawing, 2317, 2317, 4095, 4095, 0),
		(drawing, 2318, 2318, 4095, 4095, 0),
		(drawing, 2319, 2319, 4095, 4095, 0),
		(drawing, 2320, 2320, 4095, 4095, 0),
		(drawing, 2321, 2321, 4095, 4095, 0),
		(drawing, 2322, 2322, 4095, 4095, 0),
		(drawing, 2323, 2323, 4095, 4095, 0),
		(drawing, 2324, 2324, 4095, 4095, 0),
		(drawing, 2325, 2325, 4095, 4095, 0),
		(drawing, 2326, 2326, 4095, 4095, 0),
		(drawing, 2327, 2327, 4095, 4095, 0),
		(drawing, 2328, 2328, 4095, 4095, 0),
		(drawing, 2329, 2329, 4095, 4095, 0),
		(drawing, 2330, 2330, 4095, 4095, 0),
		(drawing, 2331, 2331, 4095, 4095, 0),
		(drawing, 2332, 2332, 4095, 4095, 0),
		(drawing, 2333, 2333, 4095, 4095, 0),
		(drawing, 2334, 2334, 4095, 4095, 0),
		(drawing, 2335, 2335, 4095, 4095, 0),
		(drawing, 2336, 2336, 4095, 4095, 0),
		(drawing, 2337, 2337, 4095, 4095, 0),
		(drawing, 2338, 2338, 4095, 4095, 0),
		(drawing, 2339, 2339, 4095, 4095, 0),
		(drawing, 2340, 2340, 4095, 4095, 0),
		(drawing, 2341, 2341, 4095, 4095, 0),
		(drawing, 2342, 2342, 4095, 4095, 0),
		(drawing, 2343, 2343, 4095, 4095, 0),
		(drawing, 2344, 2344, 4095, 4095, 0),
		(drawing, 2345, 2345, 4095, 4095, 0),
		(drawing, 2346, 2346, 4095, 4095, 0),
		(drawing, 2347, 2347, 4095, 4095, 0),
		(drawing, 2348, 2348, 4095, 4095, 0),
		(drawing, 2349, 2349, 4095, 4095, 0),
		(drawing, 2350, 2350, 4095, 4095, 0),
		(drawing, 2351, 2351, 4095, 4095, 0),
		(drawing, 2352, 2352, 4095, 4095, 0),
		(drawing, 2353, 2353, 4095, 4095, 0),
		(drawing, 2354, 2354, 4095, 4095, 0),
		(drawing, 2355, 2355, 4095, 4095, 0),
		(drawing, 2356, 2356, 4095, 4095, 0),
		(drawing, 2357, 2357, 4095, 4095, 0),
		(drawing, 2358, 2358, 4095, 4095, 0),
		(drawing, 2359, 2359, 4095, 4095, 0),
		(drawing, 2360, 2360, 4095, 4095, 0),
		(drawing, 2361, 2361, 4095, 4095, 0),
		(drawing, 2362, 2362, 4095, 4095, 0),
		(drawing, 2363, 2363, 4095, 4095, 0),
		(drawing, 2364, 2364, 4095, 4095, 0),
		(drawing, 2365, 2365, 4095, 4095, 0),
		(drawing, 2366, 2366, 4095, 4095, 0),
		(drawing, 2367, 2367, 4095, 4095, 0),
		(drawing, 2368, 2368, 4095, 4095, 0),
		(drawing, 2369, 2369, 4095, 4095, 0),
		(drawing, 2370, 2370, 4095, 4095, 0),
		(drawing, 2371, 2371, 4095, 4095, 0),
		(drawing, 2372, 2372, 4095, 4095, 0),
		(drawing, 2373, 2373, 4095, 4095, 0),
		(drawing, 2374, 2374, 4095, 4095, 0),
		(drawing, 2375, 2375, 4095, 4095, 0),
		(drawing, 2376, 2376, 4095, 4095, 0),
		(drawing, 2377, 2377, 4095, 4095, 0),
		(drawing, 2378, 2378, 4095, 4095, 0),
		(drawing, 2379, 2379, 4095, 4095, 0),
		(drawing, 2380, 2380, 4095, 4095, 0),
		(drawing, 2381, 2381, 4095, 4095, 0),
		(drawing, 2382, 2382, 4095, 4095, 0),
		(drawing, 2383, 2383, 4095, 4095, 0),
		(drawing, 2384, 2384, 4095, 4095, 0),
		(drawing, 2385, 2385, 4095, 4095, 0),
		(drawing, 2386, 2386, 4095, 4095, 0),
		(drawing, 2387, 2387, 4095, 4095, 0),
		(drawing, 2388, 2388, 4095, 4095, 0),
		(drawing, 2389, 2389, 4095, 4095, 0),
		(drawing, 2390, 2390, 4095, 4095, 0),
		(drawing, 2391, 2391, 4095, 4095, 0),
		(drawing, 2392, 2392, 4095, 4095, 0),
		(drawing, 2393, 2393, 4095, 4095, 0),
		(drawing, 2394, 2394, 4095, 4095, 0),
		(drawing, 2395, 2395, 4095, 4095, 0),
		(drawing, 2396, 2396, 4095, 4095, 0),
		(drawing, 2397, 2397, 4095, 4095, 0),
		(drawing, 2398, 2398, 4095, 4095, 0),
		(drawing, 2399, 2399, 4095, 4095, 0),
		(drawing, 2400, 2400, 4095, 4095, 0),
		(drawing, 2401, 2401, 4095, 4095, 0),
		(drawing, 2402, 2402, 4095, 4095, 0),
		(drawing, 2403, 2403, 4095, 4095, 0),
		(drawing, 2404, 2404, 4095, 4095, 0),
		(drawing, 2405, 2405, 4095, 4095, 0),
		(drawing, 2406, 2406, 4095, 4095, 0),
		(drawing, 2407, 2407, 4095, 4095, 0),
		(drawing, 2408, 2408, 4095, 4095, 0),
		(drawing, 2409, 2409, 4095, 4095, 0),
		(drawing, 2410, 2410, 4095, 4095, 0),
		(drawing, 2411, 2411, 4095, 4095, 0),
		(drawing, 2412, 2412, 4095, 4095, 0),
		(drawing, 2413, 2413, 4095, 4095, 0),
		(drawing, 2414, 2414, 4095, 4095, 0),
		(drawing, 2415, 2415, 4095, 4095, 0),
		(drawing, 2416, 2416, 4095, 4095, 0),
		(drawing, 2417, 2417, 4095, 4095, 0),
		(drawing, 2418, 2418, 4095, 4095, 0),
		(drawing, 2419, 2419, 4095, 4095, 0),
		(drawing, 2420, 2420, 4095, 4095, 0),
		(drawing, 2421, 2421, 4095, 4095, 0),
		(drawing, 2422, 2422, 4095, 4095, 0),
		(drawing, 2423, 2423, 4095, 4095, 0),
		(drawing, 2424, 2424, 4095, 4095, 0),
		(drawing, 2425, 2425, 4095, 4095, 0),
		(drawing, 2426, 2426, 4095, 4095, 0),
		(drawing, 2427, 2427, 4095, 4095, 0),
		(drawing, 2428, 2428, 4095, 4095, 0),
		(drawing, 2429, 2429, 4095, 4095, 0),
		(drawing, 2430, 2430, 4095, 4095, 0),
		(drawing, 2431, 2431, 4095, 4095, 0),
		(drawing, 2432, 2432, 4095, 4095, 0),
		(drawing, 2433, 2433, 4095, 4095, 0),
		(drawing, 2434, 2434, 4095, 4095, 0),
		(drawing, 2435, 2435, 4095, 4095, 0),
		(drawing, 2436, 2436, 4095, 4095, 0),
		(drawing, 2437, 2437, 4095, 4095, 0),
		(drawing, 2438, 2438, 4095, 4095, 0),
		(drawing, 2439, 2439, 4095, 4095, 0),
		(drawing, 2440, 2440, 4095, 4095, 0),
		(drawing, 2441, 2441, 4095, 4095, 0),
		(drawing, 2442, 2442, 4095, 4095, 0),
		(drawing, 2443, 2443, 4095, 4095, 0),
		(drawing, 2444, 2444, 4095, 4095, 0),
		(drawing, 2445, 2445, 4095, 4095, 0),
		(drawing, 2446, 2446, 4095, 4095, 0),
		(drawing, 2447, 2447, 4095, 4095, 0),
		(drawing, 2448, 2448, 4095, 4095, 0),
		(drawing, 2449, 2449, 4095, 4095, 0),
		(drawing, 2450, 2450, 4095, 4095, 0),
		(drawing, 2451, 2451, 4095, 4095, 0),
		(drawing, 2452, 2452, 4095, 4095, 0),
		(drawing, 2453, 2453, 4095, 4095, 0),
		(drawing, 2454, 2454, 4095, 4095, 0),
		(drawing, 2455, 2455, 4095, 4095, 0),
		(drawing, 2456, 2456, 4095, 4095, 0),
		(drawing, 2457, 2457, 4095, 4095, 0),
		(drawing, 2458, 2458, 4095, 4095, 0),
		(drawing, 2459, 2459, 4095, 4095, 0),
		(drawing, 2460, 2460, 4095, 4095, 0),
		(drawing, 2461, 2461, 4095, 4095, 0),
		(drawing, 2462, 2462, 4095, 4095, 0),
		(drawing, 2463, 2463, 4095, 4095, 0),
		(drawing, 2464, 2464, 4095, 4095, 0),
		(drawing, 2465, 2465, 4095, 4095, 0),
		(drawing, 2466, 2466, 4095, 4095, 0),
		(drawing, 2467, 2467, 4095, 4095, 0),
		(drawing, 2468, 2468, 4095, 4095, 0),
		(drawing, 2469, 2469, 4095, 4095, 0),
		(drawing, 2470, 2470, 4095, 4095, 0),
		(drawing, 2471, 2471, 4095, 4095, 0),
		(drawing, 2472, 2472, 4095, 4095, 0),
		(drawing, 2473, 2473, 4095, 4095, 0),
		(drawing, 2474, 2474, 4095, 4095, 0),
		(drawing, 2475, 2475, 4095, 4095, 0),
		(drawing, 2476, 2476, 4095, 4095, 0),
		(drawing, 2477, 2477, 4095, 4095, 0),
		(drawing, 2478, 2478, 4095, 4095, 0),
		(drawing, 2479, 2479, 4095, 4095, 0),
		(drawing, 2480, 2480, 4095, 4095, 0),
		(drawing, 2481, 2481, 4095, 4095, 0),
		(drawing, 2482, 2482, 4095, 4095, 0),
		(drawing, 2483, 2483, 4095, 4095, 0),
		(drawing, 2484, 2484, 4095, 4095, 0),
		(drawing, 2485, 2485, 4095, 4095, 0),
		(drawing, 2486, 2486, 4095, 4095, 0),
		(drawing, 2487, 2487, 4095, 4095, 0),
		(drawing, 2488, 2488, 4095, 4095, 0),
		(drawing, 2489, 2489, 4095, 4095, 0),
		(drawing, 2490, 2490, 4095, 4095, 0),
		(drawing, 2491, 2491, 4095, 4095, 0),
		(drawing, 2492, 2492, 4095, 4095, 0),
		(drawing, 2493, 2493, 4095, 4095, 0),
		(drawing, 2494, 2494, 4095, 4095, 0),
		(drawing, 2495, 2495, 4095, 4095, 0),
		(drawing, 2496, 2496, 4095, 4095, 0),
		(drawing, 2497, 2497, 4095, 4095, 0),
		(drawing, 2498, 2498, 4095, 4095, 0),
		(drawing, 2499, 2499, 4095, 4095, 0),
		(drawing, 2500, 2500, 4095, 4095, 0),
		(drawing, 2501, 2501, 4095, 4095, 0),
		(drawing, 2502, 2502, 4095, 4095, 0),
		(drawing, 2503, 2503, 4095, 4095, 0),
		(drawing, 2504, 2504, 4095, 4095, 0),
		(drawing, 2505, 2505, 4095, 4095, 0),
		(drawing, 2506, 2506, 4095, 4095, 0),
		(drawing, 2507, 2507, 4095, 4095, 0),
		(drawing, 2508, 2508, 4095, 4095, 0),
		(drawing, 2509, 2509, 4095, 4095, 0),
		(drawing, 2510, 2510, 4095, 4095, 0),
		(drawing, 2511, 2511, 4095, 4095, 0),
		(drawing, 2512, 2512, 4095, 4095, 0),
		(drawing, 2513, 2513, 4095, 4095, 0),
		(drawing, 2514, 2514, 4095, 4095, 0),
		(drawing, 2515, 2515, 4095, 4095, 0),
		(drawing, 2516, 2516, 4095, 4095, 0),
		(drawing, 2517, 2517, 4095, 4095, 0),
		(drawing, 2518, 2518, 4095, 4095, 0),
		(drawing, 2519, 2519, 4095, 4095, 0),
		(drawing, 2520, 2520, 4095, 4095, 0),
		(drawing, 2521, 2521, 4095, 4095, 0),
		(drawing, 2522, 2522, 4095, 4095, 0),
		(drawing, 2523, 2523, 4095, 4095, 0),
		(drawing, 2524, 2524, 4095, 4095, 0),
		(drawing, 2525, 2525, 4095, 4095, 0),
		(drawing, 2526, 2526, 4095, 4095, 0),
		(drawing, 2527, 2527, 4095, 4095, 0),
		(drawing, 2528, 2528, 4095, 4095, 0),
		(drawing, 2529, 2529, 4095, 4095, 0),
		(drawing, 2530, 2530, 4095, 4095, 0),
		(drawing, 2531, 2531, 4095, 4095, 0),
		(drawing, 2532, 2532, 4095, 4095, 0),
		(drawing, 2533, 2533, 4095, 4095, 0),
		(drawing, 2534, 2534, 4095, 4095, 0),
		(drawing, 2535, 2535, 4095, 4095, 0),
		(drawing, 2536, 2536, 4095, 4095, 0),
		(drawing, 2537, 2537, 4095, 4095, 0),
		(drawing, 2538, 2538, 4095, 4095, 0),
		(drawing, 2539, 2539, 4095, 4095, 0),
		(drawing, 2540, 2540, 4095, 4095, 0),
		(drawing, 2541, 2541, 4095, 4095, 0),
		(drawing, 2542, 2542, 4095, 4095, 0),
		(drawing, 2543, 2543, 4095, 4095, 0),
		(drawing, 2544, 2544, 4095, 4095, 0),
		(drawing, 2545, 2545, 4095, 4095, 0),
		(drawing, 2546, 2546, 4095, 4095, 0),
		(drawing, 2547, 2547, 4095, 4095, 0),
		(drawing, 2548, 2548, 4095, 4095, 0),
		(drawing, 2549, 2549, 4095, 4095, 0),
		(drawing, 2550, 2550, 4095, 4095, 0),
		(drawing, 2551, 2551, 4095, 4095, 0),
		(drawing, 2552, 2552, 4095, 4095, 0),
		(drawing, 2553, 2553, 4095, 4095, 0),
		(drawing, 2554, 2554, 4095, 4095, 0),
		(drawing, 2555, 2555, 4095, 4095, 0),
		(drawing, 2556, 2556, 4095, 4095, 0),
		(drawing, 2557, 2557, 4095, 4095, 0),
		(drawing, 2558, 2558, 4095, 4095, 0),
		(drawing, 2559, 2559, 4095, 4095, 0),
		(drawing, 2560, 2560, 4095, 4095, 0),
		(drawing, 2561, 2561, 4095, 4095, 0),
		(drawing, 2562, 2562, 4095, 4095, 0),
		(drawing, 2563, 2563, 4095, 4095, 0),
		(drawing, 2564, 2564, 4095, 4095, 0),
		(drawing, 2565, 2565, 4095, 4095, 0),
		(drawing, 2566, 2566, 4095, 4095, 0),
		(drawing, 2567, 2567, 4095, 4095, 0),
		(drawing, 2568, 2568, 4095, 4095, 0),
		(drawing, 2569, 2569, 4095, 4095, 0),
		(drawing, 2570, 2570, 4095, 4095, 0),
		(drawing, 2571, 2571, 4095, 4095, 0),
		(drawing, 2572, 2572, 4095, 4095, 0),
		(drawing, 2573, 2573, 4095, 4095, 0),
		(drawing, 2574, 2574, 4095, 4095, 0),
		(drawing, 2575, 2575, 4095, 4095, 0),
		(drawing, 2576, 2576, 4095, 4095, 0),
		(drawing, 2577, 2577, 4095, 4095, 0),
		(drawing, 2578, 2578, 4095, 4095, 0),
		(drawing, 2579, 2579, 4095, 4095, 0),
		(drawing, 2580, 2580, 4095, 4095, 0),
		(drawing, 2581, 2581, 4095, 4095, 0),
		(drawing, 2582, 2582, 4095, 4095, 0),
		(drawing, 2583, 2583, 4095, 4095, 0),
		(drawing, 2584, 2584, 4095, 4095, 0),
		(drawing, 2585, 2585, 4095, 4095, 0),
		(drawing, 2586, 2586, 4095, 4095, 0),
		(drawing, 2587, 2587, 4095, 4095, 0),
		(drawing, 2588, 2588, 4095, 4095, 0),
		(drawing, 2589, 2589, 4095, 4095, 0),
		(drawing, 2590, 2590, 4095, 4095, 0),
		(drawing, 2591, 2591, 4095, 4095, 0),
		(drawing, 2592, 2592, 4095, 4095, 0),
		(drawing, 2593, 2593, 4095, 4095, 0),
		(drawing, 2594, 2594, 4095, 4095, 0),
		(drawing, 2595, 2595, 4095, 4095, 0),
		(drawing, 2596, 2596, 4095, 4095, 0),
		(drawing, 2597, 2597, 4095, 4095, 0),
		(drawing, 2598, 2598, 4095, 4095, 0),
		(drawing, 2599, 2599, 4095, 4095, 0),
		(drawing, 2600, 2600, 4095, 4095, 0),
		(drawing, 2601, 2601, 4095, 4095, 0),
		(drawing, 2602, 2602, 4095, 4095, 0),
		(drawing, 2603, 2603, 4095, 4095, 0),
		(drawing, 2604, 2604, 4095, 4095, 0),
		(drawing, 2605, 2605, 4095, 4095, 0),
		(drawing, 2606, 2606, 4095, 4095, 0),
		(drawing, 2607, 2607, 4095, 4095, 0),
		(drawing, 2608, 2608, 4095, 4095, 0),
		(drawing, 2609, 2609, 4095, 4095, 0),
		(drawing, 2610, 2610, 4095, 4095, 0),
		(drawing, 2611, 2611, 4095, 4095, 0),
		(drawing, 2612, 2612, 4095, 4095, 0),
		(drawing, 2613, 2613, 4095, 4095, 0),
		(drawing, 2614, 2614, 4095, 4095, 0),
		(drawing, 2615, 2615, 4095, 4095, 0),
		(drawing, 2616, 2616, 4095, 4095, 0),
		(drawing, 2617, 2617, 4095, 4095, 0),
		(drawing, 2618, 2618, 4095, 4095, 0),
		(drawing, 2619, 2619, 4095, 4095, 0),
		(drawing, 2620, 2620, 4095, 4095, 0),
		(drawing, 2621, 2621, 4095, 4095, 0),
		(drawing, 2622, 2622, 4095, 4095, 0),
		(drawing, 2623, 2623, 4095, 4095, 0),
		(drawing, 2624, 2624, 4095, 4095, 0),
		(drawing, 2625, 2625, 4095, 4095, 0),
		(drawing, 2626, 2626, 4095, 4095, 0),
		(drawing, 2627, 2627, 4095, 4095, 0),
		(drawing, 2628, 2628, 4095, 4095, 0),
		(drawing, 2629, 2629, 4095, 4095, 0),
		(drawing, 2630, 2630, 4095, 4095, 0),
		(drawing, 2631, 2631, 4095, 4095, 0),
		(drawing, 2632, 2632, 4095, 4095, 0),
		(drawing, 2633, 2633, 4095, 4095, 0),
		(drawing, 2634, 2634, 4095, 4095, 0),
		(drawing, 2635, 2635, 4095, 4095, 0),
		(drawing, 2636, 2636, 4095, 4095, 0),
		(drawing, 2637, 2637, 4095, 4095, 0),
		(drawing, 2638, 2638, 4095, 4095, 0),
		(drawing, 2639, 2639, 4095, 4095, 0),
		(drawing, 2640, 2640, 4095, 4095, 0),
		(drawing, 2641, 2641, 4095, 4095, 0),
		(drawing, 2642, 2642, 4095, 4095, 0),
		(drawing, 2643, 2643, 4095, 4095, 0),
		(drawing, 2644, 2644, 4095, 4095, 0),
		(drawing, 2645, 2645, 4095, 4095, 0),
		(drawing, 2646, 2646, 4095, 4095, 0),
		(drawing, 2647, 2647, 4095, 4095, 0),
		(drawing, 2648, 2648, 4095, 4095, 0),
		(drawing, 2649, 2649, 4095, 4095, 0),
		(drawing, 2650, 2650, 4095, 4095, 0),
		(drawing, 2651, 2651, 4095, 4095, 0),
		(drawing, 2652, 2652, 4095, 4095, 0),
		(drawing, 2653, 2653, 4095, 4095, 0),
		(drawing, 2654, 2654, 4095, 4095, 0),
		(drawing, 2655, 2655, 4095, 4095, 0),
		(drawing, 2656, 2656, 4095, 4095, 0),
		(drawing, 2657, 2657, 4095, 4095, 0),
		(drawing, 2658, 2658, 4095, 4095, 0),
		(drawing, 2659, 2659, 4095, 4095, 0),
		(drawing, 2660, 2660, 4095, 4095, 0),
		(drawing, 2661, 2661, 4095, 4095, 0),
		(drawing, 2662, 2662, 4095, 4095, 0),
		(drawing, 2663, 2663, 4095, 4095, 0),
		(drawing, 2664, 2664, 4095, 4095, 0),
		(drawing, 2665, 2665, 4095, 4095, 0),
		(drawing, 2666, 2666, 4095, 4095, 0),
		(drawing, 2667, 2667, 4095, 4095, 0),
		(drawing, 2668, 2668, 4095, 4095, 0),
		(drawing, 2669, 2669, 4095, 4095, 0),
		(drawing, 2670, 2670, 4095, 4095, 0),
		(drawing, 2671, 2671, 4095, 4095, 0),
		(drawing, 2672, 2672, 4095, 4095, 0),
		(drawing, 2673, 2673, 4095, 4095, 0),
		(drawing, 2674, 2674, 4095, 4095, 0),
		(drawing, 2675, 2675, 4095, 4095, 0),
		(drawing, 2676, 2676, 4095, 4095, 0),
		(drawing, 2677, 2677, 4095, 4095, 0),
		(drawing, 2678, 2678, 4095, 4095, 0),
		(drawing, 2679, 2679, 4095, 4095, 0),
		(drawing, 2680, 2680, 4095, 4095, 0),
		(drawing, 2681, 2681, 4095, 4095, 0),
		(drawing, 2682, 2682, 4095, 4095, 0),
		(drawing, 2683, 2683, 4095, 4095, 0),
		(drawing, 2684, 2684, 4095, 4095, 0),
		(drawing, 2685, 2685, 4095, 4095, 0),
		(drawing, 2686, 2686, 4095, 4095, 0),
		(drawing, 2687, 2687, 4095, 4095, 0),
		(drawing, 2688, 2688, 4095, 4095, 0),
		(drawing, 2689, 2689, 4095, 4095, 0),
		(drawing, 2690, 2690, 4095, 4095, 0),
		(drawing, 2691, 2691, 4095, 4095, 0),
		(drawing, 2692, 2692, 4095, 4095, 0),
		(drawing, 2693, 2693, 4095, 4095, 0),
		(drawing, 2694, 2694, 4095, 4095, 0),
		(drawing, 2695, 2695, 4095, 4095, 0),
		(drawing, 2696, 2696, 4095, 4095, 0),
		(drawing, 2697, 2697, 4095, 4095, 0),
		(drawing, 2698, 2698, 4095, 4095, 0),
		(drawing, 2699, 2699, 4095, 4095, 0),
		(drawing, 2700, 2700, 4095, 4095, 0),
		(drawing, 2701, 2701, 4095, 4095, 0),
		(drawing, 2702, 2702, 4095, 4095, 0),
		(drawing, 2703, 2703, 4095, 4095, 0),
		(drawing, 2704, 2704, 4095, 4095, 0),
		(drawing, 2705, 2705, 4095, 4095, 0),
		(drawing, 2706, 2706, 4095, 4095, 0),
		(drawing, 2707, 2707, 4095, 4095, 0),
		(drawing, 2708, 2708, 4095, 4095, 0),
		(drawing, 2709, 2709, 4095, 4095, 0),
		(drawing, 2710, 2710, 4095, 4095, 0),
		(drawing, 2711, 2711, 4095, 4095, 0),
		(drawing, 2712, 2712, 4095, 4095, 0),
		(drawing, 2713, 2713, 4095, 4095, 0),
		(drawing, 2714, 2714, 4095, 4095, 0),
		(drawing, 2715, 2715, 4095, 4095, 0),
		(drawing, 2716, 2716, 4095, 4095, 0),
		(drawing, 2717, 2717, 4095, 4095, 0),
		(drawing, 2718, 2718, 4095, 4095, 0),
		(drawing, 2719, 2719, 4095, 4095, 0),
		(drawing, 2720, 2720, 4095, 4095, 0),
		(drawing, 2721, 2721, 4095, 4095, 0),
		(drawing, 2722, 2722, 4095, 4095, 0),
		(drawing, 2723, 2723, 4095, 4095, 0),
		(drawing, 2724, 2724, 4095, 4095, 0),
		(drawing, 2725, 2725, 4095, 4095, 0),
		(drawing, 2726, 2726, 4095, 4095, 0),
		(drawing, 2727, 2727, 4095, 4095, 0),
		(drawing, 2728, 2728, 4095, 4095, 0),
		(drawing, 2729, 2729, 4095, 4095, 0),
		(drawing, 2730, 2730, 4095, 4095, 0),
		(drawing, 2731, 2731, 4095, 4095, 0),
		(drawing, 2732, 2732, 4095, 4095, 0),
		(drawing, 2733, 2733, 4095, 4095, 0),
		(drawing, 2734, 2734, 4095, 4095, 0),
		(drawing, 2735, 2735, 4095, 4095, 0),
		(drawing, 2736, 2736, 4095, 4095, 0),
		(drawing, 2737, 2737, 4095, 4095, 0),
		(drawing, 2738, 2738, 4095, 4095, 0),
		(drawing, 2739, 2739, 4095, 4095, 0),
		(drawing, 2740, 2740, 4095, 4095, 0),
		(drawing, 2741, 2741, 4095, 4095, 0),
		(drawing, 2742, 2742, 4095, 4095, 0),
		(drawing, 2743, 2743, 4095, 4095, 0),
		(drawing, 2744, 2744, 4095, 4095, 0),
		(drawing, 2745, 2745, 4095, 4095, 0),
		(drawing, 2746, 2746, 4095, 4095, 0),
		(drawing, 2747, 2747, 4095, 4095, 0),
		(drawing, 2748, 2748, 4095, 4095, 0),
		(drawing, 2749, 2749, 4095, 4095, 0),
		(drawing, 2750, 2750, 4095, 4095, 0),
		(drawing, 2751, 2751, 4095, 4095, 0),
		(drawing, 2752, 2752, 4095, 4095, 0),
		(drawing, 2753, 2753, 4095, 4095, 0),
		(drawing, 2754, 2754, 4095, 4095, 0),
		(drawing, 2755, 2755, 4095, 4095, 0),
		(drawing, 2756, 2756, 4095, 4095, 0),
		(drawing, 2757, 2757, 4095, 4095, 0),
		(drawing, 2758, 2758, 4095, 4095, 0),
		(drawing, 2759, 2759, 4095, 4095, 0),
		(drawing, 2760, 2760, 4095, 4095, 0),
		(drawing, 2761, 2761, 4095, 4095, 0),
		(drawing, 2762, 2762, 4095, 4095, 0),
		(drawing, 2763, 2763, 4095, 4095, 0),
		(drawing, 2764, 2764, 4095, 4095, 0),
		(drawing, 2765, 2765, 4095, 4095, 0),
		(drawing, 2766, 2766, 4095, 4095, 0),
		(drawing, 2767, 2767, 4095, 4095, 0),
		(drawing, 2768, 2768, 4095, 4095, 0),
		(drawing, 2769, 2769, 4095, 4095, 0),
		(drawing, 2770, 2770, 4095, 4095, 0),
		(drawing, 2771, 2771, 4095, 4095, 0),
		(drawing, 2772, 2772, 4095, 4095, 0),
		(drawing, 2773, 2773, 4095, 4095, 0),
		(drawing, 2774, 2774, 4095, 4095, 0),
		(drawing, 2775, 2775, 4095, 4095, 0),
		(drawing, 2776, 2776, 4095, 4095, 0),
		(drawing, 2777, 2777, 4095, 4095, 0),
		(drawing, 2778, 2778, 4095, 4095, 0),
		(drawing, 2779, 2779, 4095, 4095, 0),
		(drawing, 2780, 2780, 4095, 4095, 0),
		(drawing, 2781, 2781, 4095, 4095, 0),
		(drawing, 2782, 2782, 4095, 4095, 0),
		(drawing, 2783, 2783, 4095, 4095, 0),
		(drawing, 2784, 2784, 4095, 4095, 0),
		(drawing, 2785, 2785, 4095, 4095, 0),
		(drawing, 2786, 2786, 4095, 4095, 0),
		(drawing, 2787, 2787, 4095, 4095, 0),
		(drawing, 2788, 2788, 4095, 4095, 0),
		(drawing, 2789, 2789, 4095, 4095, 0),
		(drawing, 2790, 2790, 4095, 4095, 0),
		(drawing, 2791, 2791, 4095, 4095, 0),
		(drawing, 2792, 2792, 4095, 4095, 0),
		(drawing, 2793, 2793, 4095, 4095, 0),
		(drawing, 2794, 2794, 4095, 4095, 0),
		(drawing, 2795, 2795, 4095, 4095, 0),
		(drawing, 2796, 2796, 4095, 4095, 0),
		(drawing, 2797, 2797, 4095, 4095, 0),
		(drawing, 2798, 2798, 4095, 4095, 0),
		(drawing, 2799, 2799, 4095, 4095, 0),
		(drawing, 2800, 2800, 4095, 4095, 0),
		(drawing, 2801, 2801, 4095, 4095, 0),
		(drawing, 2802, 2802, 4095, 4095, 0),
		(drawing, 2803, 2803, 4095, 4095, 0),
		(drawing, 2804, 2804, 4095, 4095, 0),
		(drawing, 2805, 2805, 4095, 4095, 0),
		(drawing, 2806, 2806, 4095, 4095, 0),
		(drawing, 2807, 2807, 4095, 4095, 0),
		(drawing, 2808, 2808, 4095, 4095, 0),
		(drawing, 2809, 2809, 4095, 4095, 0),
		(drawing, 2810, 2810, 4095, 4095, 0),
		(drawing, 2811, 2811, 4095, 4095, 0),
		(drawing, 2812, 2812, 4095, 4095, 0),
		(drawing, 2813, 2813, 4095, 4095, 0),
		(drawing, 2814, 2814, 4095, 4095, 0),
		(drawing, 2815, 2815, 4095, 4095, 0),
		(drawing, 2816, 2816, 4095, 4095, 0),
		(drawing, 2817, 2817, 4095, 4095, 0),
		(drawing, 2818, 2818, 4095, 4095, 0),
		(drawing, 2819, 2819, 4095, 4095, 0),
		(drawing, 2820, 2820, 4095, 4095, 0),
		(drawing, 2821, 2821, 4095, 4095, 0),
		(drawing, 2822, 2822, 4095, 4095, 0),
		(drawing, 2823, 2823, 4095, 4095, 0),
		(drawing, 2824, 2824, 4095, 4095, 0),
		(drawing, 2825, 2825, 4095, 4095, 0),
		(drawing, 2826, 2826, 4095, 4095, 0),
		(drawing, 2827, 2827, 4095, 4095, 0),
		(drawing, 2828, 2828, 4095, 4095, 0),
		(drawing, 2829, 2829, 4095, 4095, 0),
		(drawing, 2830, 2830, 4095, 4095, 0),
		(drawing, 2831, 2831, 4095, 4095, 0),
		(drawing, 2832, 2832, 4095, 4095, 0),
		(drawing, 2833, 2833, 4095, 4095, 0),
		(drawing, 2834, 2834, 4095, 4095, 0),
		(drawing, 2835, 2835, 4095, 4095, 0),
		(drawing, 2836, 2836, 4095, 4095, 0),
		(drawing, 2837, 2837, 4095, 4095, 0),
		(drawing, 2838, 2838, 4095, 4095, 0),
		(drawing, 2839, 2839, 4095, 4095, 0),
		(drawing, 2840, 2840, 4095, 4095, 0),
		(drawing, 2841, 2841, 4095, 4095, 0),
		(drawing, 2842, 2842, 4095, 4095, 0),
		(drawing, 2843, 2843, 4095, 4095, 0),
		(drawing, 2844, 2844, 4095, 4095, 0),
		(drawing, 2845, 2845, 4095, 4095, 0),
		(drawing, 2846, 2846, 4095, 4095, 0),
		(drawing, 2847, 2847, 4095, 4095, 0),
		(drawing, 2848, 2848, 4095, 4095, 0),
		(drawing, 2849, 2849, 4095, 4095, 0),
		(drawing, 2850, 2850, 4095, 4095, 0),
		(drawing, 2851, 2851, 4095, 4095, 0),
		(drawing, 2852, 2852, 4095, 4095, 0),
		(drawing, 2853, 2853, 4095, 4095, 0),
		(drawing, 2854, 2854, 4095, 4095, 0),
		(drawing, 2855, 2855, 4095, 4095, 0),
		(drawing, 2856, 2856, 4095, 4095, 0),
		(drawing, 2857, 2857, 4095, 4095, 0),
		(drawing, 2858, 2858, 4095, 4095, 0),
		(drawing, 2859, 2859, 4095, 4095, 0),
		(drawing, 2860, 2860, 4095, 4095, 0),
		(drawing, 2861, 2861, 4095, 4095, 0),
		(drawing, 2862, 2862, 4095, 4095, 0),
		(drawing, 2863, 2863, 4095, 4095, 0),
		(drawing, 2864, 2864, 4095, 4095, 0),
		(drawing, 2865, 2865, 4095, 4095, 0),
		(drawing, 2866, 2866, 4095, 4095, 0),
		(drawing, 2867, 2867, 4095, 4095, 0),
		(drawing, 2868, 2868, 4095, 4095, 0),
		(drawing, 2869, 2869, 4095, 4095, 0),
		(drawing, 2870, 2870, 4095, 4095, 0),
		(drawing, 2871, 2871, 4095, 4095, 0),
		(drawing, 2872, 2872, 4095, 4095, 0),
		(drawing, 2873, 2873, 4095, 4095, 0),
		(drawing, 2874, 2874, 4095, 4095, 0),
		(drawing, 2875, 2875, 4095, 4095, 0),
		(drawing, 2876, 2876, 4095, 4095, 0),
		(drawing, 2877, 2877, 4095, 4095, 0),
		(drawing, 2878, 2878, 4095, 4095, 0),
		(drawing, 2879, 2879, 4095, 4095, 0),
		(drawing, 2880, 2880, 4095, 4095, 0),
		(drawing, 2881, 2881, 4095, 4095, 0),
		(drawing, 2882, 2882, 4095, 4095, 0),
		(drawing, 2883, 2883, 4095, 4095, 0),
		(drawing, 2884, 2884, 4095, 4095, 0),
		(drawing, 2885, 2885, 4095, 4095, 0),
		(drawing, 2886, 2886, 4095, 4095, 0),
		(drawing, 2887, 2887, 4095, 4095, 0),
		(drawing, 2888, 2888, 4095, 4095, 0),
		(drawing, 2889, 2889, 4095, 4095, 0),
		(drawing, 2890, 2890, 4095, 4095, 0),
		(drawing, 2891, 2891, 4095, 4095, 0),
		(drawing, 2892, 2892, 4095, 4095, 0),
		(drawing, 2893, 2893, 4095, 4095, 0),
		(drawing, 2894, 2894, 4095, 4095, 0),
		(drawing, 2895, 2895, 4095, 4095, 0),
		(drawing, 2896, 2896, 4095, 4095, 0),
		(drawing, 2897, 2897, 4095, 4095, 0),
		(drawing, 2898, 2898, 4095, 4095, 0),
		(drawing, 2899, 2899, 4095, 4095, 0),
		(drawing, 2900, 2900, 4095, 4095, 0),
		(drawing, 2901, 2901, 4095, 4095, 0),
		(drawing, 2902, 2902, 4095, 4095, 0),
		(drawing, 2903, 2903, 4095, 4095, 0),
		(drawing, 2904, 2904, 4095, 4095, 0),
		(drawing, 2905, 2905, 4095, 4095, 0),
		(drawing, 2906, 2906, 4095, 4095, 0),
		(drawing, 2907, 2907, 4095, 4095, 0),
		(drawing, 2908, 2908, 4095, 4095, 0),
		(drawing, 2909, 2909, 4095, 4095, 0),
		(drawing, 2910, 2910, 4095, 4095, 0),
		(drawing, 2911, 2911, 4095, 4095, 0),
		(drawing, 2912, 2912, 4095, 4095, 0),
		(drawing, 2913, 2913, 4095, 4095, 0),
		(drawing, 2914, 2914, 4095, 4095, 0),
		(drawing, 2915, 2915, 4095, 4095, 0),
		(drawing, 2916, 2916, 4095, 4095, 0),
		(drawing, 2917, 2917, 4095, 4095, 0),
		(drawing, 2918, 2918, 4095, 4095, 0),
		(drawing, 2919, 2919, 4095, 4095, 0),
		(drawing, 2920, 2920, 4095, 4095, 0),
		(drawing, 2921, 2921, 4095, 4095, 0),
		(drawing, 2922, 2922, 4095, 4095, 0),
		(drawing, 2923, 2923, 4095, 4095, 0),
		(drawing, 2924, 2924, 4095, 4095, 0),
		(drawing, 2925, 2925, 4095, 4095, 0),
		(drawing, 2926, 2926, 4095, 4095, 0),
		(drawing, 2927, 2927, 4095, 4095, 0),
		(drawing, 2928, 2928, 4095, 4095, 0),
		(drawing, 2929, 2929, 4095, 4095, 0),
		(drawing, 2930, 2930, 4095, 4095, 0),
		(drawing, 2931, 2931, 4095, 4095, 0),
		(drawing, 2932, 2932, 4095, 4095, 0),
		(drawing, 2933, 2933, 4095, 4095, 0),
		(drawing, 2934, 2934, 4095, 4095, 0),
		(drawing, 2935, 2935, 4095, 4095, 0),
		(drawing, 2936, 2936, 4095, 4095, 0),
		(drawing, 2937, 2937, 4095, 4095, 0),
		(drawing, 2938, 2938, 4095, 4095, 0),
		(drawing, 2939, 2939, 4095, 4095, 0),
		(drawing, 2940, 2940, 4095, 4095, 0),
		(drawing, 2941, 2941, 4095, 4095, 0),
		(drawing, 2942, 2942, 4095, 4095, 0),
		(drawing, 2943, 2943, 4095, 4095, 0),
		(drawing, 2944, 2944, 4095, 4095, 0),
		(drawing, 2945, 2945, 4095, 4095, 0),
		(drawing, 2946, 2946, 4095, 4095, 0),
		(drawing, 2947, 2947, 4095, 4095, 0),
		(drawing, 2948, 2948, 4095, 4095, 0),
		(drawing, 2949, 2949, 4095, 4095, 0),
		(drawing, 2950, 2950, 4095, 4095, 0),
		(drawing, 2951, 2951, 4095, 4095, 0),
		(drawing, 2952, 2952, 4095, 4095, 0),
		(drawing, 2953, 2953, 4095, 4095, 0),
		(drawing, 2954, 2954, 4095, 4095, 0),
		(drawing, 2955, 2955, 4095, 4095, 0),
		(drawing, 2956, 2956, 4095, 4095, 0),
		(drawing, 2957, 2957, 4095, 4095, 0),
		(drawing, 2958, 2958, 4095, 4095, 0),
		(drawing, 2959, 2959, 4095, 4095, 0),
		(drawing, 2960, 2960, 4095, 4095, 0),
		(drawing, 2961, 2961, 4095, 4095, 0),
		(drawing, 2962, 2962, 4095, 4095, 0),
		(drawing, 2963, 2963, 4095, 4095, 0),
		(drawing, 2964, 2964, 4095, 4095, 0),
		(drawing, 2965, 2965, 4095, 4095, 0),
		(drawing, 2966, 2966, 4095, 4095, 0),
		(drawing, 2967, 2967, 4095, 4095, 0),
		(drawing, 2968, 2968, 4095, 4095, 0),
		(drawing, 2969, 2969, 4095, 4095, 0),
		(drawing, 2970, 2970, 4095, 4095, 0),
		(drawing, 2971, 2971, 4095, 4095, 0),
		(drawing, 2972, 2972, 4095, 4095, 0),
		(drawing, 2973, 2973, 4095, 4095, 0),
		(drawing, 2974, 2974, 4095, 4095, 0),
		(drawing, 2975, 2975, 4095, 4095, 0),
		(drawing, 2976, 2976, 4095, 4095, 0),
		(drawing, 2977, 2977, 4095, 4095, 0),
		(drawing, 2978, 2978, 4095, 4095, 0),
		(drawing, 2979, 2979, 4095, 4095, 0),
		(drawing, 2980, 2980, 4095, 4095, 0),
		(drawing, 2981, 2981, 4095, 4095, 0),
		(drawing, 2982, 2982, 4095, 4095, 0),
		(drawing, 2983, 2983, 4095, 4095, 0),
		(drawing, 2984, 2984, 4095, 4095, 0),
		(drawing, 2985, 2985, 4095, 4095, 0),
		(drawing, 2986, 2986, 4095, 4095, 0),
		(drawing, 2987, 2987, 4095, 4095, 0),
		(drawing, 2988, 2988, 4095, 4095, 0),
		(drawing, 2989, 2989, 4095, 4095, 0),
		(drawing, 2990, 2990, 4095, 4095, 0),
		(drawing, 2991, 2991, 4095, 4095, 0),
		(drawing, 2992, 2992, 4095, 4095, 0),
		(drawing, 2993, 2993, 4095, 4095, 0),
		(drawing, 2994, 2994, 4095, 4095, 0),
		(drawing, 2995, 2995, 4095, 4095, 0),
		(drawing, 2996, 2996, 4095, 4095, 0),
		(drawing, 2997, 2997, 4095, 4095, 0),
		(drawing, 2998, 2998, 4095, 4095, 0),
		(drawing, 2999, 2999, 4095, 4095, 0),
		(drawing, 3000, 3000, 4095, 4095, 0),
		(drawing, 3001, 3001, 4095, 4095, 0),
		(drawing, 3002, 3002, 4095, 4095, 0),
		(drawing, 3003, 3003, 4095, 4095, 0),
		(drawing, 3004, 3004, 4095, 4095, 0),
		(drawing, 3005, 3005, 4095, 4095, 0),
		(drawing, 3006, 3006, 4095, 4095, 0),
		(drawing, 3007, 3007, 4095, 4095, 0),
		(drawing, 3008, 3008, 4095, 4095, 0),
		(drawing, 3009, 3009, 4095, 4095, 0),
		(drawing, 3010, 3010, 4095, 4095, 0),
		(drawing, 3011, 3011, 4095, 4095, 0),
		(drawing, 3012, 3012, 4095, 4095, 0),
		(drawing, 3013, 3013, 4095, 4095, 0),
		(drawing, 3014, 3014, 4095, 4095, 0),
		(drawing, 3015, 3015, 4095, 4095, 0),
		(drawing, 3016, 3016, 4095, 4095, 0),
		(drawing, 3017, 3017, 4095, 4095, 0),
		(drawing, 3018, 3018, 4095, 4095, 0),
		(drawing, 3019, 3019, 4095, 4095, 0),
		(drawing, 3020, 3020, 4095, 4095, 0),
		(drawing, 3021, 3021, 4095, 4095, 0),
		(drawing, 3022, 3022, 4095, 4095, 0),
		(drawing, 3023, 3023, 4095, 4095, 0),
		(drawing, 3024, 3024, 4095, 4095, 0),
		(drawing, 3025, 3025, 4095, 4095, 0),
		(drawing, 3026, 3026, 4095, 4095, 0),
		(drawing, 3027, 3027, 4095, 4095, 0),
		(drawing, 3028, 3028, 4095, 4095, 0),
		(drawing, 3029, 3029, 4095, 4095, 0),
		(drawing, 3030, 3030, 4095, 4095, 0),
		(drawing, 3031, 3031, 4095, 4095, 0),
		(drawing, 3032, 3032, 4095, 4095, 0),
		(drawing, 3033, 3033, 4095, 4095, 0),
		(drawing, 3034, 3034, 4095, 4095, 0),
		(drawing, 3035, 3035, 4095, 4095, 0),
		(drawing, 3036, 3036, 4095, 4095, 0),
		(drawing, 3037, 3037, 4095, 4095, 0),
		(drawing, 3038, 3038, 4095, 4095, 0),
		(drawing, 3039, 3039, 4095, 4095, 0),
		(drawing, 3040, 3040, 4095, 4095, 0),
		(drawing, 3041, 3041, 4095, 4095, 0),
		(drawing, 3042, 3042, 4095, 4095, 0),
		(drawing, 3043, 3043, 4095, 4095, 0),
		(drawing, 3044, 3044, 4095, 4095, 0),
		(drawing, 3045, 3045, 4095, 4095, 0),
		(drawing, 3046, 3046, 4095, 4095, 0),
		(drawing, 3047, 3047, 4095, 4095, 0),
		(drawing, 3048, 3048, 4095, 4095, 0),
		(drawing, 3049, 3049, 4095, 4095, 0),
		(drawing, 3050, 3050, 4095, 4095, 0),
		(drawing, 3051, 3051, 4095, 4095, 0),
		(drawing, 3052, 3052, 4095, 4095, 0),
		(drawing, 3053, 3053, 4095, 4095, 0),
		(drawing, 3054, 3054, 4095, 4095, 0),
		(drawing, 3055, 3055, 4095, 4095, 0),
		(drawing, 3056, 3056, 4095, 4095, 0),
		(drawing, 3057, 3057, 4095, 4095, 0),
		(drawing, 3058, 3058, 4095, 4095, 0),
		(drawing, 3059, 3059, 4095, 4095, 0),
		(drawing, 3060, 3060, 4095, 4095, 0),
		(drawing, 3061, 3061, 4095, 4095, 0),
		(drawing, 3062, 3062, 4095, 4095, 0),
		(drawing, 3063, 3063, 4095, 4095, 0),
		(drawing, 3064, 3064, 4095, 4095, 0),
		(drawing, 3065, 3065, 4095, 4095, 0),
		(drawing, 3066, 3066, 4095, 4095, 0),
		(drawing, 3067, 3067, 4095, 4095, 0),
		(drawing, 3068, 3068, 4095, 4095, 0),
		(drawing, 3069, 3069, 4095, 4095, 0),
		(drawing, 3070, 3070, 4095, 4095, 0),
		(drawing, 3071, 3071, 4095, 4095, 0),
		(drawing, 3072, 3072, 4095, 4095, 0),
		(drawing, 3073, 3073, 4095, 4095, 0),
		(drawing, 3074, 3074, 4095, 4095, 0),
		(drawing, 3075, 3075, 4095, 4095, 0),
		(drawing, 3076, 3076, 4095, 4095, 0),
		(drawing, 3077, 3077, 4095, 4095, 0),
		(drawing, 3078, 3078, 4095, 4095, 0),
		(drawing, 3079, 3079, 4095, 4095, 0),
		(drawing, 3080, 3080, 4095, 4095, 0),
		(drawing, 3081, 3081, 4095, 4095, 0),
		(drawing, 3082, 3082, 4095, 4095, 0),
		(drawing, 3083, 3083, 4095, 4095, 0),
		(drawing, 3084, 3084, 4095, 4095, 0),
		(drawing, 3085, 3085, 4095, 4095, 0),
		(drawing, 3086, 3086, 4095, 4095, 0),
		(drawing, 3087, 3087, 4095, 4095, 0),
		(drawing, 3088, 3088, 4095, 4095, 0),
		(drawing, 3089, 3089, 4095, 4095, 0),
		(drawing, 3090, 3090, 4095, 4095, 0),
		(drawing, 3091, 3091, 4095, 4095, 0),
		(drawing, 3092, 3092, 4095, 4095, 0),
		(drawing, 3093, 3093, 4095, 4095, 0),
		(drawing, 3094, 3094, 4095, 4095, 0),
		(drawing, 3095, 3095, 4095, 4095, 0),
		(drawing, 3096, 3096, 4095, 4095, 0),
		(drawing, 3097, 3097, 4095, 4095, 0),
		(drawing, 3098, 3098, 4095, 4095, 0),
		(drawing, 3099, 3099, 4095, 4095, 0),
		(drawing, 3100, 3100, 4095, 4095, 0),
		(drawing, 3101, 3101, 4095, 4095, 0),
		(drawing, 3102, 3102, 4095, 4095, 0),
		(drawing, 3103, 3103, 4095, 4095, 0),
		(drawing, 3104, 3104, 4095, 4095, 0),
		(drawing, 3105, 3105, 4095, 4095, 0),
		(drawing, 3106, 3106, 4095, 4095, 0),
		(drawing, 3107, 3107, 4095, 4095, 0),
		(drawing, 3108, 3108, 4095, 4095, 0),
		(drawing, 3109, 3109, 4095, 4095, 0),
		(drawing, 3110, 3110, 4095, 4095, 0),
		(drawing, 3111, 3111, 4095, 4095, 0),
		(drawing, 3112, 3112, 4095, 4095, 0),
		(drawing, 3113, 3113, 4095, 4095, 0),
		(drawing, 3114, 3114, 4095, 4095, 0),
		(drawing, 3115, 3115, 4095, 4095, 0),
		(drawing, 3116, 3116, 4095, 4095, 0),
		(drawing, 3117, 3117, 4095, 4095, 0),
		(drawing, 3118, 3118, 4095, 4095, 0),
		(drawing, 3119, 3119, 4095, 4095, 0),
		(drawing, 3120, 3120, 4095, 4095, 0),
		(drawing, 3121, 3121, 4095, 4095, 0),
		(drawing, 3122, 3122, 4095, 4095, 0),
		(drawing, 3123, 3123, 4095, 4095, 0),
		(drawing, 3124, 3124, 4095, 4095, 0),
		(drawing, 3125, 3125, 4095, 4095, 0),
		(drawing, 3126, 3126, 4095, 4095, 0),
		(drawing, 3127, 3127, 4095, 4095, 0),
		(drawing, 3128, 3128, 4095, 4095, 0),
		(drawing, 3129, 3129, 4095, 4095, 0),
		(drawing, 3130, 3130, 4095, 4095, 0),
		(drawing, 3131, 3131, 4095, 4095, 0),
		(drawing, 3132, 3132, 4095, 4095, 0),
		(drawing, 3133, 3133, 4095, 4095, 0),
		(drawing, 3134, 3134, 4095, 4095, 0),
		(drawing, 3135, 3135, 4095, 4095, 0),
		(drawing, 3136, 3136, 4095, 4095, 0),
		(drawing, 3137, 3137, 4095, 4095, 0),
		(drawing, 3138, 3138, 4095, 4095, 0),
		(drawing, 3139, 3139, 4095, 4095, 0),
		(drawing, 3140, 3140, 4095, 4095, 0),
		(drawing, 3141, 3141, 4095, 4095, 0),
		(drawing, 3142, 3142, 4095, 4095, 0),
		(drawing, 3143, 3143, 4095, 4095, 0),
		(drawing, 3144, 3144, 4095, 4095, 0),
		(drawing, 3145, 3145, 4095, 4095, 0),
		(drawing, 3146, 3146, 4095, 4095, 0),
		(drawing, 3147, 3147, 4095, 4095, 0),
		(drawing, 3148, 3148, 4095, 4095, 0),
		(drawing, 3149, 3149, 4095, 4095, 0),
		(drawing, 3150, 3150, 4095, 4095, 0),
		(drawing, 3151, 3151, 4095, 4095, 0),
		(drawing, 3152, 3152, 4095, 4095, 0),
		(drawing, 3153, 3153, 4095, 4095, 0),
		(drawing, 3154, 3154, 4095, 4095, 0),
		(drawing, 3155, 3155, 4095, 4095, 0),
		(drawing, 3156, 3156, 4095, 4095, 0),
		(drawing, 3157, 3157, 4095, 4095, 0),
		(drawing, 3158, 3158, 4095, 4095, 0),
		(drawing, 3159, 3159, 4095, 4095, 0),
		(drawing, 3160, 3160, 4095, 4095, 0),
		(drawing, 3161, 3161, 4095, 4095, 0),
		(drawing, 3162, 3162, 4095, 4095, 0),
		(drawing, 3163, 3163, 4095, 4095, 0),
		(drawing, 3164, 3164, 4095, 4095, 0),
		(drawing, 3165, 3165, 4095, 4095, 0),
		(drawing, 3166, 3166, 4095, 4095, 0),
		(drawing, 3167, 3167, 4095, 4095, 0),
		(drawing, 3168, 3168, 4095, 4095, 0),
		(drawing, 3169, 3169, 4095, 4095, 0),
		(drawing, 3170, 3170, 4095, 4095, 0),
		(drawing, 3171, 3171, 4095, 4095, 0),
		(drawing, 3172, 3172, 4095, 4095, 0),
		(drawing, 3173, 3173, 4095, 4095, 0),
		(drawing, 3174, 3174, 4095, 4095, 0),
		(drawing, 3175, 3175, 4095, 4095, 0),
		(drawing, 3176, 3176, 4095, 4095, 0),
		(drawing, 3177, 3177, 4095, 4095, 0),
		(drawing, 3178, 3178, 4095, 4095, 0),
		(drawing, 3179, 3179, 4095, 4095, 0),
		(drawing, 3180, 3180, 4095, 4095, 0),
		(drawing, 3181, 3181, 4095, 4095, 0),
		(drawing, 3182, 3182, 4095, 4095, 0),
		(drawing, 3183, 3183, 4095, 4095, 0),
		(drawing, 3184, 3184, 4095, 4095, 0),
		(drawing, 3185, 3185, 4095, 4095, 0),
		(drawing, 3186, 3186, 4095, 4095, 0),
		(drawing, 3187, 3187, 4095, 4095, 0),
		(drawing, 3188, 3188, 4095, 4095, 0),
		(drawing, 3189, 3189, 4095, 4095, 0),
		(drawing, 3190, 3190, 4095, 4095, 0),
		(drawing, 3191, 3191, 4095, 4095, 0),
		(drawing, 3192, 3192, 4095, 4095, 0),
		(drawing, 3193, 3193, 4095, 4095, 0),
		(drawing, 3194, 3194, 4095, 4095, 0),
		(drawing, 3195, 3195, 4095, 4095, 0),
		(drawing, 3196, 3196, 4095, 4095, 0),
		(drawing, 3197, 3197, 4095, 4095, 0),
		(drawing, 3198, 3198, 4095, 4095, 0),
		(drawing, 3199, 3199, 4095, 4095, 0),
		(drawing, 3200, 3200, 4095, 4095, 0),
		(drawing, 3201, 3201, 4095, 4095, 0),
		(drawing, 3202, 3202, 4095, 4095, 0),
		(drawing, 3203, 3203, 4095, 4095, 0),
		(drawing, 3204, 3204, 4095, 4095, 0),
		(drawing, 3205, 3205, 4095, 4095, 0),
		(drawing, 3206, 3206, 4095, 4095, 0),
		(drawing, 3207, 3207, 4095, 4095, 0),
		(drawing, 3208, 3208, 4095, 4095, 0),
		(drawing, 3209, 3209, 4095, 4095, 0),
		(drawing, 3210, 3210, 4095, 4095, 0),
		(drawing, 3211, 3211, 4095, 4095, 0),
		(drawing, 3212, 3212, 4095, 4095, 0),
		(drawing, 3213, 3213, 4095, 4095, 0),
		(drawing, 3214, 3214, 4095, 4095, 0),
		(drawing, 3215, 3215, 4095, 4095, 0),
		(drawing, 3216, 3216, 4095, 4095, 0),
		(drawing, 3217, 3217, 4095, 4095, 0),
		(drawing, 3218, 3218, 4095, 4095, 0),
		(drawing, 3219, 3219, 4095, 4095, 0),
		(drawing, 3220, 3220, 4095, 4095, 0),
		(drawing, 3221, 3221, 4095, 4095, 0),
		(drawing, 3222, 3222, 4095, 4095, 0),
		(drawing, 3223, 3223, 4095, 4095, 0),
		(drawing, 3224, 3224, 4095, 4095, 0),
		(drawing, 3225, 3225, 4095, 4095, 0),
		(drawing, 3226, 3226, 4095, 4095, 0),
		(drawing, 3227, 3227, 4095, 4095, 0),
		(drawing, 3228, 3228, 4095, 4095, 0),
		(drawing, 3229, 3229, 4095, 4095, 0),
		(drawing, 3230, 3230, 4095, 4095, 0),
		(drawing, 3231, 3231, 4095, 4095, 0),
		(drawing, 3232, 3232, 4095, 4095, 0),
		(drawing, 3233, 3233, 4095, 4095, 0),
		(drawing, 3234, 3234, 4095, 4095, 0),
		(drawing, 3235, 3235, 4095, 4095, 0),
		(drawing, 3236, 3236, 4095, 4095, 0),
		(drawing, 3237, 3237, 4095, 4095, 0),
		(drawing, 3238, 3238, 4095, 4095, 0),
		(drawing, 3239, 3239, 4095, 4095, 0),
		(drawing, 3240, 3240, 4095, 4095, 0),
		(drawing, 3241, 3241, 4095, 4095, 0),
		(drawing, 3242, 3242, 4095, 4095, 0),
		(drawing, 3243, 3243, 4095, 4095, 0),
		(drawing, 3244, 3244, 4095, 4095, 0),
		(drawing, 3245, 3245, 4095, 4095, 0),
		(drawing, 3246, 3246, 4095, 4095, 0),
		(drawing, 3247, 3247, 4095, 4095, 0),
		(drawing, 3248, 3248, 4095, 4095, 0),
		(drawing, 3249, 3249, 4095, 4095, 0),
		(drawing, 3250, 3250, 4095, 4095, 0),
		(drawing, 3251, 3251, 4095, 4095, 0),
		(drawing, 3252, 3252, 4095, 4095, 0),
		(drawing, 3253, 3253, 4095, 4095, 0),
		(drawing, 3254, 3254, 4095, 4095, 0),
		(drawing, 3255, 3255, 4095, 4095, 0),
		(drawing, 3256, 3256, 4095, 4095, 0),
		(drawing, 3257, 3257, 4095, 4095, 0),
		(drawing, 3258, 3258, 4095, 4095, 0),
		(drawing, 3259, 3259, 4095, 4095, 0),
		(drawing, 3260, 3260, 4095, 4095, 0),
		(drawing, 3261, 3261, 4095, 4095, 0),
		(drawing, 3262, 3262, 4095, 4095, 0),
		(drawing, 3263, 3263, 4095, 4095, 0),
		(drawing, 3264, 3264, 4095, 4095, 0),
		(drawing, 3265, 3265, 4095, 4095, 0),
		(drawing, 3266, 3266, 4095, 4095, 0),
		(drawing, 3267, 3267, 4095, 4095, 0),
		(drawing, 3268, 3268, 4095, 4095, 0),
		(drawing, 3269, 3269, 4095, 4095, 0),
		(drawing, 3270, 3270, 4095, 4095, 0),
		(drawing, 3271, 3271, 4095, 4095, 0),
		(drawing, 3272, 3272, 4095, 4095, 0),
		(drawing, 3273, 3273, 4095, 4095, 0),
		(drawing, 3274, 3274, 4095, 4095, 0),
		(drawing, 3275, 3275, 4095, 4095, 0),
		(drawing, 3276, 3276, 4095, 4095, 0),
		(drawing, 3277, 3277, 4095, 4095, 0),
		(drawing, 3278, 3278, 4095, 4095, 0),
		(drawing, 3279, 3279, 4095, 4095, 0),
		(drawing, 3280, 3280, 4095, 4095, 0),
		(drawing, 3281, 3281, 4095, 4095, 0),
		(drawing, 3282, 3282, 4095, 4095, 0),
		(drawing, 3283, 3283, 4095, 4095, 0),
		(drawing, 3284, 3284, 4095, 4095, 0),
		(drawing, 3285, 3285, 4095, 4095, 0),
		(drawing, 3286, 3286, 4095, 4095, 0),
		(drawing, 3287, 3287, 4095, 4095, 0),
		(drawing, 3288, 3288, 4095, 4095, 0),
		(drawing, 3289, 3289, 4095, 4095, 0),
		(drawing, 3290, 3290, 4095, 4095, 0),
		(drawing, 3291, 3291, 4095, 4095, 0),
		(drawing, 3292, 3292, 4095, 4095, 0),
		(drawing, 3293, 3293, 4095, 4095, 0),
		(drawing, 3294, 3294, 4095, 4095, 0),
		(drawing, 3295, 3295, 4095, 4095, 0),
		(drawing, 3296, 3296, 4095, 4095, 0),
		(drawing, 3297, 3297, 4095, 4095, 0),
		(drawing, 3298, 3298, 4095, 4095, 0),
		(drawing, 3299, 3299, 4095, 4095, 0),
		(drawing, 3300, 3300, 4095, 4095, 0),
		(drawing, 3301, 3301, 4095, 4095, 0),
		(drawing, 3302, 3302, 4095, 4095, 0),
		(drawing, 3303, 3303, 4095, 4095, 0),
		(drawing, 3304, 3304, 4095, 4095, 0),
		(drawing, 3305, 3305, 4095, 4095, 0),
		(drawing, 3306, 3306, 4095, 4095, 0),
		(drawing, 3307, 3307, 4095, 4095, 0),
		(drawing, 3308, 3308, 4095, 4095, 0),
		(drawing, 3309, 3309, 4095, 4095, 0),
		(drawing, 3310, 3310, 4095, 4095, 0),
		(drawing, 3311, 3311, 4095, 4095, 0),
		(drawing, 3312, 3312, 4095, 4095, 0),
		(drawing, 3313, 3313, 4095, 4095, 0),
		(drawing, 3314, 3314, 4095, 4095, 0),
		(drawing, 3315, 3315, 4095, 4095, 0),
		(drawing, 3316, 3316, 4095, 4095, 0),
		(drawing, 3317, 3317, 4095, 4095, 0),
		(drawing, 3318, 3318, 4095, 4095, 0),
		(drawing, 3319, 3319, 4095, 4095, 0),
		(drawing, 3320, 3320, 4095, 4095, 0),
		(drawing, 3321, 3321, 4095, 4095, 0),
		(drawing, 3322, 3322, 4095, 4095, 0),
		(drawing, 3323, 3323, 4095, 4095, 0),
		(drawing, 3324, 3324, 4095, 4095, 0),
		(drawing, 3325, 3325, 4095, 4095, 0),
		(drawing, 3326, 3326, 4095, 4095, 0),
		(drawing, 3327, 3327, 4095, 4095, 0),
		(drawing, 3328, 3328, 4095, 4095, 0),
		(drawing, 3329, 3329, 4095, 4095, 0),
		(drawing, 3330, 3330, 4095, 4095, 0),
		(drawing, 3331, 3331, 4095, 4095, 0),
		(drawing, 3332, 3332, 4095, 4095, 0),
		(drawing, 3333, 3333, 4095, 4095, 0),
		(drawing, 3334, 3334, 4095, 4095, 0),
		(drawing, 3335, 3335, 4095, 4095, 0),
		(drawing, 3336, 3336, 4095, 4095, 0),
		(drawing, 3337, 3337, 4095, 4095, 0),
		(drawing, 3338, 3338, 4095, 4095, 0),
		(drawing, 3339, 3339, 4095, 4095, 0),
		(drawing, 3340, 3340, 4095, 4095, 0),
		(drawing, 3341, 3341, 4095, 4095, 0),
		(drawing, 3342, 3342, 4095, 4095, 0),
		(drawing, 3343, 3343, 4095, 4095, 0),
		(drawing, 3344, 3344, 4095, 4095, 0),
		(drawing, 3345, 3345, 4095, 4095, 0),
		(drawing, 3346, 3346, 4095, 4095, 0),
		(drawing, 3347, 3347, 4095, 4095, 0),
		(drawing, 3348, 3348, 4095, 4095, 0),
		(drawing, 3349, 3349, 4095, 4095, 0),
		(drawing, 3350, 3350, 4095, 4095, 0),
		(drawing, 3351, 3351, 4095, 4095, 0),
		(drawing, 3352, 3352, 4095, 4095, 0),
		(drawing, 3353, 3353, 4095, 4095, 0),
		(drawing, 3354, 3354, 4095, 4095, 0),
		(drawing, 3355, 3355, 4095, 4095, 0),
		(drawing, 3356, 3356, 4095, 4095, 0),
		(drawing, 3357, 3357, 4095, 4095, 0),
		(drawing, 3358, 3358, 4095, 4095, 0),
		(drawing, 3359, 3359, 4095, 4095, 0),
		(drawing, 3360, 3360, 4095, 4095, 0),
		(drawing, 3361, 3361, 4095, 4095, 0),
		(drawing, 3362, 3362, 4095, 4095, 0),
		(drawing, 3363, 3363, 4095, 4095, 0),
		(drawing, 3364, 3364, 4095, 4095, 0),
		(drawing, 3365, 3365, 4095, 4095, 0),
		(drawing, 3366, 3366, 4095, 4095, 0),
		(drawing, 3367, 3367, 4095, 4095, 0),
		(drawing, 3368, 3368, 4095, 4095, 0),
		(drawing, 3369, 3369, 4095, 4095, 0),
		(drawing, 3370, 3370, 4095, 4095, 0),
		(drawing, 3371, 3371, 4095, 4095, 0),
		(drawing, 3372, 3372, 4095, 4095, 0),
		(drawing, 3373, 3373, 4095, 4095, 0),
		(drawing, 3374, 3374, 4095, 4095, 0),
		(drawing, 3375, 3375, 4095, 4095, 0),
		(drawing, 3376, 3376, 4095, 4095, 0),
		(drawing, 3377, 3377, 4095, 4095, 0),
		(drawing, 3378, 3378, 4095, 4095, 0),
		(drawing, 3379, 3379, 4095, 4095, 0),
		(drawing, 3380, 3380, 4095, 4095, 0),
		(drawing, 3381, 3381, 4095, 4095, 0),
		(drawing, 3382, 3382, 4095, 4095, 0),
		(drawing, 3383, 3383, 4095, 4095, 0),
		(drawing, 3384, 3384, 4095, 4095, 0),
		(drawing, 3385, 3385, 4095, 4095, 0),
		(drawing, 3386, 3386, 4095, 4095, 0),
		(drawing, 3387, 3387, 4095, 4095, 0),
		(drawing, 3388, 3388, 4095, 4095, 0),
		(drawing, 3389, 3389, 4095, 4095, 0),
		(drawing, 3390, 3390, 4095, 4095, 0),
		(drawing, 3391, 3391, 4095, 4095, 0),
		(drawing, 3392, 3392, 4095, 4095, 0),
		(drawing, 3393, 3393, 4095, 4095, 0),
		(drawing, 3394, 3394, 4095, 4095, 0),
		(drawing, 3395, 3395, 4095, 4095, 0),
		(drawing, 3396, 3396, 4095, 4095, 0),
		(drawing, 3397, 3397, 4095, 4095, 0),
		(drawing, 3398, 3398, 4095, 4095, 0),
		(drawing, 3399, 3399, 4095, 4095, 0),
		(drawing, 3400, 3400, 4095, 4095, 0),
		(drawing, 3401, 3401, 4095, 4095, 0),
		(drawing, 3402, 3402, 4095, 4095, 0),
		(drawing, 3403, 3403, 4095, 4095, 0),
		(drawing, 3404, 3404, 4095, 4095, 0),
		(drawing, 3405, 3405, 4095, 4095, 0),
		(drawing, 3406, 3406, 4095, 4095, 0),
		(drawing, 3407, 3407, 4095, 4095, 0),
		(drawing, 3408, 3408, 4095, 4095, 0),
		(drawing, 3409, 3409, 4095, 4095, 0),
		(drawing, 3410, 3410, 4095, 4095, 0),
		(drawing, 3411, 3411, 4095, 4095, 0),
		(drawing, 3412, 3412, 4095, 4095, 0),
		(drawing, 3413, 3413, 4095, 4095, 0),
		(drawing, 3414, 3414, 4095, 4095, 0),
		(drawing, 3415, 3415, 4095, 4095, 0),
		(drawing, 3416, 3416, 4095, 4095, 0),
		(drawing, 3417, 3417, 4095, 4095, 0),
		(drawing, 3418, 3418, 4095, 4095, 0),
		(drawing, 3419, 3419, 4095, 4095, 0),
		(drawing, 3420, 3420, 4095, 4095, 0),
		(drawing, 3421, 3421, 4095, 4095, 0),
		(drawing, 3422, 3422, 4095, 4095, 0),
		(drawing, 3423, 3423, 4095, 4095, 0),
		(drawing, 3424, 3424, 4095, 4095, 0),
		(drawing, 3425, 3425, 4095, 4095, 0),
		(drawing, 3426, 3426, 4095, 4095, 0),
		(drawing, 3427, 3427, 4095, 4095, 0),
		(drawing, 3428, 3428, 4095, 4095, 0),
		(drawing, 3429, 3429, 4095, 4095, 0),
		(drawing, 3430, 3430, 4095, 4095, 0),
		(drawing, 3431, 3431, 4095, 4095, 0),
		(drawing, 3432, 3432, 4095, 4095, 0),
		(drawing, 3433, 3433, 4095, 4095, 0),
		(drawing, 3434, 3434, 4095, 4095, 0),
		(drawing, 3435, 3435, 4095, 4095, 0),
		(drawing, 3436, 3436, 4095, 4095, 0),
		(drawing, 3437, 3437, 4095, 4095, 0),
		(drawing, 3438, 3438, 4095, 4095, 0),
		(drawing, 3439, 3439, 4095, 4095, 0),
		(drawing, 3440, 3440, 4095, 4095, 0),
		(drawing, 3441, 3441, 4095, 4095, 0),
		(drawing, 3442, 3442, 4095, 4095, 0),
		(drawing, 3443, 3443, 4095, 4095, 0),
		(drawing, 3444, 3444, 4095, 4095, 0),
		(drawing, 3445, 3445, 4095, 4095, 0),
		(drawing, 3446, 3446, 4095, 4095, 0),
		(drawing, 3447, 3447, 4095, 4095, 0),
		(drawing, 3448, 3448, 4095, 4095, 0),
		(drawing, 3449, 3449, 4095, 4095, 0),
		(drawing, 3450, 3450, 4095, 4095, 0),
		(drawing, 3451, 3451, 4095, 4095, 0),
		(drawing, 3452, 3452, 4095, 4095, 0),
		(drawing, 3453, 3453, 4095, 4095, 0),
		(drawing, 3454, 3454, 4095, 4095, 0),
		(drawing, 3455, 3455, 4095, 4095, 0),
		(drawing, 3456, 3456, 4095, 4095, 0),
		(drawing, 3457, 3457, 4095, 4095, 0),
		(drawing, 3458, 3458, 4095, 4095, 0),
		(drawing, 3459, 3459, 4095, 4095, 0),
		(drawing, 3460, 3460, 4095, 4095, 0),
		(drawing, 3461, 3461, 4095, 4095, 0),
		(drawing, 3462, 3462, 4095, 4095, 0),
		(drawing, 3463, 3463, 4095, 4095, 0),
		(drawing, 3464, 3464, 4095, 4095, 0),
		(drawing, 3465, 3465, 4095, 4095, 0),
		(drawing, 3466, 3466, 4095, 4095, 0),
		(drawing, 3467, 3467, 4095, 4095, 0),
		(drawing, 3468, 3468, 4095, 4095, 0),
		(drawing, 3469, 3469, 4095, 4095, 0),
		(drawing, 3470, 3470, 4095, 4095, 0),
		(drawing, 3471, 3471, 4095, 4095, 0),
		(drawing, 3472, 3472, 4095, 4095, 0),
		(drawing, 3473, 3473, 4095, 4095, 0),
		(drawing, 3474, 3474, 4095, 4095, 0),
		(drawing, 3475, 3475, 4095, 4095, 0),
		(drawing, 3476, 3476, 4095, 4095, 0),
		(drawing, 3477, 3477, 4095, 4095, 0),
		(drawing, 3478, 3478, 4095, 4095, 0),
		(drawing, 3479, 3479, 4095, 4095, 0),
		(drawing, 3480, 3480, 4095, 4095, 0),
		(drawing, 3481, 3481, 4095, 4095, 0),
		(drawing, 3482, 3482, 4095, 4095, 0),
		(drawing, 3483, 3483, 4095, 4095, 0),
		(drawing, 3484, 3484, 4095, 4095, 0),
		(drawing, 3485, 3485, 4095, 4095, 0),
		(drawing, 3486, 3486, 4095, 4095, 0),
		(drawing, 3487, 3487, 4095, 4095, 0),
		(drawing, 3488, 3488, 4095, 4095, 0),
		(drawing, 3489, 3489, 4095, 4095, 0),
		(drawing, 3490, 3490, 4095, 4095, 0),
		(drawing, 3491, 3491, 4095, 4095, 0),
		(drawing, 3492, 3492, 4095, 4095, 0),
		(drawing, 3493, 3493, 4095, 4095, 0),
		(drawing, 3494, 3494, 4095, 4095, 0),
		(drawing, 3495, 3495, 4095, 4095, 0),
		(drawing, 3496, 3496, 4095, 4095, 0),
		(drawing, 3497, 3497, 4095, 4095, 0),
		(drawing, 3498, 3498, 4095, 4095, 0),
		(drawing, 3499, 3499, 4095, 4095, 0),
		(drawing, 3500, 3500, 4095, 4095, 0),
		(drawing, 3501, 3501, 4095, 4095, 0),
		(drawing, 3502, 3502, 4095, 4095, 0),
		(drawing, 3503, 3503, 4095, 4095, 0),
		(drawing, 3504, 3504, 4095, 4095, 0),
		(drawing, 3505, 3505, 4095, 4095, 0),
		(drawing, 3506, 3506, 4095, 4095, 0),
		(drawing, 3507, 3507, 4095, 4095, 0),
		(drawing, 3508, 3508, 4095, 4095, 0),
		(drawing, 3509, 3509, 4095, 4095, 0),
		(drawing, 3510, 3510, 4095, 4095, 0),
		(drawing, 3511, 3511, 4095, 4095, 0),
		(drawing, 3512, 3512, 4095, 4095, 0),
		(drawing, 3513, 3513, 4095, 4095, 0),
		(drawing, 3514, 3514, 4095, 4095, 0),
		(drawing, 3515, 3515, 4095, 4095, 0),
		(drawing, 3516, 3516, 4095, 4095, 0),
		(drawing, 3517, 3517, 4095, 4095, 0),
		(drawing, 3518, 3518, 4095, 4095, 0),
		(drawing, 3519, 3519, 4095, 4095, 0),
		(drawing, 3520, 3520, 4095, 4095, 0),
		(drawing, 3521, 3521, 4095, 4095, 0),
		(drawing, 3522, 3522, 4095, 4095, 0),
		(drawing, 3523, 3523, 4095, 4095, 0),
		(drawing, 3524, 3524, 4095, 4095, 0),
		(drawing, 3525, 3525, 4095, 4095, 0),
		(drawing, 3526, 3526, 4095, 4095, 0),
		(drawing, 3527, 3527, 4095, 4095, 0),
		(drawing, 3528, 3528, 4095, 4095, 0),
		(drawing, 3529, 3529, 4095, 4095, 0),
		(drawing, 3530, 3530, 4095, 4095, 0),
		(drawing, 3531, 3531, 4095, 4095, 0),
		(drawing, 3532, 3532, 4095, 4095, 0),
		(drawing, 3533, 3533, 4095, 4095, 0),
		(drawing, 3534, 3534, 4095, 4095, 0),
		(drawing, 3535, 3535, 4095, 4095, 0),
		(drawing, 3536, 3536, 4095, 4095, 0),
		(drawing, 3537, 3537, 4095, 4095, 0),
		(drawing, 3538, 3538, 4095, 4095, 0),
		(drawing, 3539, 3539, 4095, 4095, 0),
		(drawing, 3540, 3540, 4095, 4095, 0),
		(drawing, 3541, 3541, 4095, 4095, 0),
		(drawing, 3542, 3542, 4095, 4095, 0),
		(drawing, 3543, 3543, 4095, 4095, 0),
		(drawing, 3544, 3544, 4095, 4095, 0),
		(drawing, 3545, 3545, 4095, 4095, 0),
		(drawing, 3546, 3546, 4095, 4095, 0),
		(drawing, 3547, 3547, 4095, 4095, 0),
		(drawing, 3548, 3548, 4095, 4095, 0),
		(drawing, 3549, 3549, 4095, 4095, 0),
		(drawing, 3550, 3550, 4095, 4095, 0),
		(drawing, 3551, 3551, 4095, 4095, 0),
		(drawing, 3552, 3552, 4095, 4095, 0),
		(drawing, 3553, 3553, 4095, 4095, 0),
		(drawing, 3554, 3554, 4095, 4095, 0),
		(drawing, 3555, 3555, 4095, 4095, 0),
		(drawing, 3556, 3556, 4095, 4095, 0),
		(drawing, 3557, 3557, 4095, 4095, 0),
		(drawing, 3558, 3558, 4095, 4095, 0),
		(drawing, 3559, 3559, 4095, 4095, 0),
		(drawing, 3560, 3560, 4095, 4095, 0),
		(drawing, 3561, 3561, 4095, 4095, 0),
		(drawing, 3562, 3562, 4095, 4095, 0),
		(drawing, 3563, 3563, 4095, 4095, 0),
		(drawing, 3564, 3564, 4095, 4095, 0),
		(drawing, 3565, 3565, 4095, 4095, 0),
		(drawing, 3566, 3566, 4095, 4095, 0),
		(drawing, 3567, 3567, 4095, 4095, 0),
		(drawing, 3568, 3568, 4095, 4095, 0),
		(drawing, 3569, 3569, 4095, 4095, 0),
		(drawing, 3570, 3570, 4095, 4095, 0),
		(drawing, 3571, 3571, 4095, 4095, 0),
		(drawing, 3572, 3572, 4095, 4095, 0),
		(drawing, 3573, 3573, 4095, 4095, 0),
		(drawing, 3574, 3574, 4095, 4095, 0),
		(drawing, 3575, 3575, 4095, 4095, 0),
		(drawing, 3576, 3576, 4095, 4095, 0),
		(drawing, 3577, 3577, 4095, 4095, 0),
		(drawing, 3578, 3578, 4095, 4095, 0),
		(drawing, 3579, 3579, 4095, 4095, 0),
		(drawing, 3580, 3580, 4095, 4095, 0),
		(drawing, 3581, 3581, 4095, 4095, 0),
		(drawing, 3582, 3582, 4095, 4095, 0),
		(drawing, 3583, 3583, 4095, 4095, 0),
		(drawing, 3584, 3584, 4095, 4095, 0),
		(drawing, 3585, 3585, 4095, 4095, 0),
		(drawing, 3586, 3586, 4095, 4095, 0),
		(drawing, 3587, 3587, 4095, 4095, 0),
		(drawing, 3588, 3588, 4095, 4095, 0),
		(drawing, 3589, 3589, 4095, 4095, 0),
		(drawing, 3590, 3590, 4095, 4095, 0),
		(drawing, 3591, 3591, 4095, 4095, 0),
		(drawing, 3592, 3592, 4095, 4095, 0),
		(drawing, 3593, 3593, 4095, 4095, 0),
		(drawing, 3594, 3594, 4095, 4095, 0),
		(drawing, 3595, 3595, 4095, 4095, 0),
		(drawing, 3596, 3596, 4095, 4095, 0),
		(drawing, 3597, 3597, 4095, 4095, 0),
		(drawing, 3598, 3598, 4095, 4095, 0),
		(drawing, 3599, 3599, 4095, 4095, 0),
		(drawing, 3600, 3600, 4095, 4095, 0),
		(drawing, 3601, 3601, 4095, 4095, 0),
		(drawing, 3602, 3602, 4095, 4095, 0),
		(drawing, 3603, 3603, 4095, 4095, 0),
		(drawing, 3604, 3604, 4095, 4095, 0),
		(drawing, 3605, 3605, 4095, 4095, 0),
		(drawing, 3606, 3606, 4095, 4095, 0),
		(drawing, 3607, 3607, 4095, 4095, 0),
		(drawing, 3608, 3608, 4095, 4095, 0),
		(drawing, 3609, 3609, 4095, 4095, 0),
		(drawing, 3610, 3610, 4095, 4095, 0),
		(drawing, 3611, 3611, 4095, 4095, 0),
		(drawing, 3612, 3612, 4095, 4095, 0),
		(drawing, 3613, 3613, 4095, 4095, 0),
		(drawing, 3614, 3614, 4095, 4095, 0),
		(drawing, 3615, 3615, 4095, 4095, 0),
		(drawing, 3616, 3616, 4095, 4095, 0),
		(drawing, 3617, 3617, 4095, 4095, 0),
		(drawing, 3618, 3618, 4095, 4095, 0),
		(drawing, 3619, 3619, 4095, 4095, 0),
		(drawing, 3620, 3620, 4095, 4095, 0),
		(drawing, 3621, 3621, 4095, 4095, 0),
		(drawing, 3622, 3622, 4095, 4095, 0),
		(drawing, 3623, 3623, 4095, 4095, 0),
		(drawing, 3624, 3624, 4095, 4095, 0),
		(drawing, 3625, 3625, 4095, 4095, 0),
		(drawing, 3626, 3626, 4095, 4095, 0),
		(drawing, 3627, 3627, 4095, 4095, 0),
		(drawing, 3628, 3628, 4095, 4095, 0),
		(drawing, 3629, 3629, 4095, 4095, 0),
		(drawing, 3630, 3630, 4095, 4095, 0),
		(drawing, 3631, 3631, 4095, 4095, 0),
		(drawing, 3632, 3632, 4095, 4095, 0),
		(drawing, 3633, 3633, 4095, 4095, 0),
		(drawing, 3634, 3634, 4095, 4095, 0),
		(drawing, 3635, 3635, 4095, 4095, 0),
		(drawing, 3636, 3636, 4095, 4095, 0),
		(drawing, 3637, 3637, 4095, 4095, 0),
		(drawing, 3638, 3638, 4095, 4095, 0),
		(drawing, 3639, 3639, 4095, 4095, 0),
		(drawing, 3640, 3640, 4095, 4095, 0),
		(drawing, 3641, 3641, 4095, 4095, 0),
		(drawing, 3642, 3642, 4095, 4095, 0),
		(drawing, 3643, 3643, 4095, 4095, 0),
		(drawing, 3644, 3644, 4095, 4095, 0),
		(drawing, 3645, 3645, 4095, 4095, 0),
		(drawing, 3646, 3646, 4095, 4095, 0),
		(drawing, 3647, 3647, 4095, 4095, 0),
		(drawing, 3648, 3648, 4095, 4095, 0),
		(drawing, 3649, 3649, 4095, 4095, 0),
		(drawing, 3650, 3650, 4095, 4095, 0),
		(drawing, 3651, 3651, 4095, 4095, 0),
		(drawing, 3652, 3652, 4095, 4095, 0),
		(drawing, 3653, 3653, 4095, 4095, 0),
		(drawing, 3654, 3654, 4095, 4095, 0),
		(drawing, 3655, 3655, 4095, 4095, 0),
		(drawing, 3656, 3656, 4095, 4095, 0),
		(drawing, 3657, 3657, 4095, 4095, 0),
		(drawing, 3658, 3658, 4095, 4095, 0),
		(drawing, 3659, 3659, 4095, 4095, 0),
		(drawing, 3660, 3660, 4095, 4095, 0),
		(drawing, 3661, 3661, 4095, 4095, 0),
		(drawing, 3662, 3662, 4095, 4095, 0),
		(drawing, 3663, 3663, 4095, 4095, 0),
		(drawing, 3664, 3664, 4095, 4095, 0),
		(drawing, 3665, 3665, 4095, 4095, 0),
		(drawing, 3666, 3666, 4095, 4095, 0),
		(drawing, 3667, 3667, 4095, 4095, 0),
		(drawing, 3668, 3668, 4095, 4095, 0),
		(drawing, 3669, 3669, 4095, 4095, 0),
		(drawing, 3670, 3670, 4095, 4095, 0),
		(drawing, 3671, 3671, 4095, 4095, 0),
		(drawing, 3672, 3672, 4095, 4095, 0),
		(drawing, 3673, 3673, 4095, 4095, 0),
		(drawing, 3674, 3674, 4095, 4095, 0),
		(drawing, 3675, 3675, 4095, 4095, 0),
		(drawing, 3676, 3676, 4095, 4095, 0),
		(drawing, 3677, 3677, 4095, 4095, 0),
		(drawing, 3678, 3678, 4095, 4095, 0),
		(drawing, 3679, 3679, 4095, 4095, 0),
		(drawing, 3680, 3680, 4095, 4095, 0),
		(drawing, 3681, 3681, 4095, 4095, 0),
		(drawing, 3682, 3682, 4095, 4095, 0),
		(drawing, 3683, 3683, 4095, 4095, 0),
		(drawing, 3684, 3684, 4095, 4095, 0),
		(drawing, 3685, 3685, 4095, 4095, 0),
		(drawing, 3686, 3686, 4095, 4095, 0),
		(drawing, 3687, 3687, 4095, 4095, 0),
		(drawing, 3688, 3688, 4095, 4095, 0),
		(drawing, 3689, 3689, 4095, 4095, 0),
		(drawing, 3690, 3690, 4095, 4095, 0),
		(drawing, 3691, 3691, 4095, 4095, 0),
		(drawing, 3692, 3692, 4095, 4095, 0),
		(drawing, 3693, 3693, 4095, 4095, 0),
		(drawing, 3694, 3694, 4095, 4095, 0),
		(drawing, 3695, 3695, 4095, 4095, 0),
		(drawing, 3696, 3696, 4095, 4095, 0),
		(drawing, 3697, 3697, 4095, 4095, 0),
		(drawing, 3698, 3698, 4095, 4095, 0),
		(drawing, 3699, 3699, 4095, 4095, 0),
		(drawing, 3700, 3700, 4095, 4095, 0),
		(drawing, 3701, 3701, 4095, 4095, 0),
		(drawing, 3702, 3702, 4095, 4095, 0),
		(drawing, 3703, 3703, 4095, 4095, 0),
		(drawing, 3704, 3704, 4095, 4095, 0),
		(drawing, 3705, 3705, 4095, 4095, 0),
		(drawing, 3706, 3706, 4095, 4095, 0),
		(drawing, 3707, 3707, 4095, 4095, 0),
		(drawing, 3708, 3708, 4095, 4095, 0),
		(drawing, 3709, 3709, 4095, 4095, 0),
		(drawing, 3710, 3710, 4095, 4095, 0),
		(drawing, 3711, 3711, 4095, 4095, 0),
		(drawing, 3712, 3712, 4095, 4095, 0),
		(drawing, 3713, 3713, 4095, 4095, 0),
		(drawing, 3714, 3714, 4095, 4095, 0),
		(drawing, 3715, 3715, 4095, 4095, 0),
		(drawing, 3716, 3716, 4095, 4095, 0),
		(drawing, 3717, 3717, 4095, 4095, 0),
		(drawing, 3718, 3718, 4095, 4095, 0),
		(drawing, 3719, 3719, 4095, 4095, 0),
		(drawing, 3720, 3720, 4095, 4095, 0),
		(drawing, 3721, 3721, 4095, 4095, 0),
		(drawing, 3722, 3722, 4095, 4095, 0),
		(drawing, 3723, 3723, 4095, 4095, 0),
		(drawing, 3724, 3724, 4095, 4095, 0),
		(drawing, 3725, 3725, 4095, 4095, 0),
		(drawing, 3726, 3726, 4095, 4095, 0),
		(drawing, 3727, 3727, 4095, 4095, 0),
		(drawing, 3728, 3728, 4095, 4095, 0),
		(drawing, 3729, 3729, 4095, 4095, 0),
		(drawing, 3730, 3730, 4095, 4095, 0),
		(drawing, 3731, 3731, 4095, 4095, 0),
		(drawing, 3732, 3732, 4095, 4095, 0),
		(drawing, 3733, 3733, 4095, 4095, 0),
		(drawing, 3734, 3734, 4095, 4095, 0),
		(drawing, 3735, 3735, 4095, 4095, 0),
		(drawing, 3736, 3736, 4095, 4095, 0),
		(drawing, 3737, 3737, 4095, 4095, 0),
		(drawing, 3738, 3738, 4095, 4095, 0),
		(drawing, 3739, 3739, 4095, 4095, 0),
		(drawing, 3740, 3740, 4095, 4095, 0),
		(drawing, 3741, 3741, 4095, 4095, 0),
		(drawing, 3742, 3742, 4095, 4095, 0),
		(drawing, 3743, 3743, 4095, 4095, 0),
		(drawing, 3744, 3744, 4095, 4095, 0),
		(drawing, 3745, 3745, 4095, 4095, 0),
		(drawing, 3746, 3746, 4095, 4095, 0),
		(drawing, 3747, 3747, 4095, 4095, 0),
		(drawing, 3748, 3748, 4095, 4095, 0),
		(drawing, 3749, 3749, 4095, 4095, 0),
		(drawing, 3750, 3750, 4095, 4095, 0),
		(drawing, 3751, 3751, 4095, 4095, 0),
		(drawing, 3752, 3752, 4095, 4095, 0),
		(drawing, 3753, 3753, 4095, 4095, 0),
		(drawing, 3754, 3754, 4095, 4095, 0),
		(drawing, 3755, 3755, 4095, 4095, 0),
		(drawing, 3756, 3756, 4095, 4095, 0),
		(drawing, 3757, 3757, 4095, 4095, 0),
		(drawing, 3758, 3758, 4095, 4095, 0),
		(drawing, 3759, 3759, 4095, 4095, 0),
		(drawing, 3760, 3760, 4095, 4095, 0),
		(drawing, 3761, 3761, 4095, 4095, 0),
		(drawing, 3762, 3762, 4095, 4095, 0),
		(drawing, 3763, 3763, 4095, 4095, 0),
		(drawing, 3764, 3764, 4095, 4095, 0),
		(drawing, 3765, 3765, 4095, 4095, 0),
		(drawing, 3766, 3766, 4095, 4095, 0),
		(drawing, 3767, 3767, 4095, 4095, 0),
		(drawing, 3768, 3768, 4095, 4095, 0),
		(drawing, 3769, 3769, 4095, 4095, 0),
		(drawing, 3770, 3770, 4095, 4095, 0),
		(drawing, 3771, 3771, 4095, 4095, 0),
		(drawing, 3772, 3772, 4095, 4095, 0),
		(drawing, 3773, 3773, 4095, 4095, 0),
		(drawing, 3774, 3774, 4095, 4095, 0),
		(drawing, 3775, 3775, 4095, 4095, 0),
		(drawing, 3776, 3776, 4095, 4095, 0),
		(drawing, 3777, 3777, 4095, 4095, 0),
		(drawing, 3778, 3778, 4095, 4095, 0),
		(drawing, 3779, 3779, 4095, 4095, 0),
		(drawing, 3780, 3780, 4095, 4095, 0),
		(drawing, 3781, 3781, 4095, 4095, 0),
		(drawing, 3782, 3782, 4095, 4095, 0),
		(drawing, 3783, 3783, 4095, 4095, 0),
		(drawing, 3784, 3784, 4095, 4095, 0),
		(drawing, 3785, 3785, 4095, 4095, 0),
		(drawing, 3786, 3786, 4095, 4095, 0),
		(drawing, 3787, 3787, 4095, 4095, 0),
		(drawing, 3788, 3788, 4095, 4095, 0),
		(drawing, 3789, 3789, 4095, 4095, 0),
		(drawing, 3790, 3790, 4095, 4095, 0),
		(drawing, 3791, 3791, 4095, 4095, 0),
		(drawing, 3792, 3792, 4095, 4095, 0),
		(drawing, 3793, 3793, 4095, 4095, 0),
		(drawing, 3794, 3794, 4095, 4095, 0),
		(drawing, 3795, 3795, 4095, 4095, 0),
		(drawing, 3796, 3796, 4095, 4095, 0),
		(drawing, 3797, 3797, 4095, 4095, 0),
		(drawing, 3798, 3798, 4095, 4095, 0),
		(drawing, 3799, 3799, 4095, 4095, 0),
		(drawing, 3800, 3800, 4095, 4095, 0),
		(drawing, 3801, 3801, 4095, 4095, 0),
		(drawing, 3802, 3802, 4095, 4095, 0),
		(drawing, 3803, 3803, 4095, 4095, 0),
		(drawing, 3804, 3804, 4095, 4095, 0),
		(drawing, 3805, 3805, 4095, 4095, 0),
		(drawing, 3806, 3806, 4095, 4095, 0),
		(drawing, 3807, 3807, 4095, 4095, 0),
		(drawing, 3808, 3808, 4095, 4095, 0),
		(drawing, 3809, 3809, 4095, 4095, 0),
		(drawing, 3810, 3810, 4095, 4095, 0),
		(drawing, 3811, 3811, 4095, 4095, 0),
		(drawing, 3812, 3812, 4095, 4095, 0),
		(drawing, 3813, 3813, 4095, 4095, 0),
		(drawing, 3814, 3814, 4095, 4095, 0),
		(drawing, 3815, 3815, 4095, 4095, 0),
		(drawing, 3816, 3816, 4095, 4095, 0),
		(drawing, 3817, 3817, 4095, 4095, 0),
		(drawing, 3818, 3818, 4095, 4095, 0),
		(drawing, 3819, 3819, 4095, 4095, 0),
		(drawing, 3820, 3820, 4095, 4095, 0),
		(drawing, 3821, 3821, 4095, 4095, 0),
		(drawing, 3822, 3822, 4095, 4095, 0),
		(drawing, 3823, 3823, 4095, 4095, 0),
		(drawing, 3824, 3824, 4095, 4095, 0),
		(drawing, 3825, 3825, 4095, 4095, 0),
		(drawing, 3826, 3826, 4095, 4095, 0),
		(drawing, 3827, 3827, 4095, 4095, 0),
		(drawing, 3828, 3828, 4095, 4095, 0),
		(drawing, 3829, 3829, 4095, 4095, 0),
		(drawing, 3830, 3830, 4095, 4095, 0),
		(drawing, 3831, 3831, 4095, 4095, 0),
		(drawing, 3832, 3832, 4095, 4095, 0),
		(drawing, 3833, 3833, 4095, 4095, 0),
		(drawing, 3834, 3834, 4095, 4095, 0),
		(drawing, 3835, 3835, 4095, 4095, 0),
		(drawing, 3836, 3836, 4095, 4095, 0),
		(drawing, 3837, 3837, 4095, 4095, 0),
		(drawing, 3838, 3838, 4095, 4095, 0),
		(drawing, 3839, 3839, 4095, 4095, 0),
		(drawing, 3840, 3840, 4095, 4095, 0),
		(drawing, 3841, 3841, 4095, 4095, 0),
		(drawing, 3842, 3842, 4095, 4095, 0),
		(drawing, 3843, 3843, 4095, 4095, 0),
		(drawing, 3844, 3844, 4095, 4095, 0),
		(drawing, 3845, 3845, 4095, 4095, 0),
		(drawing, 3846, 3846, 4095, 4095, 0),
		(drawing, 3847, 3847, 4095, 4095, 0),
		(drawing, 3848, 3848, 4095, 4095, 0),
		(drawing, 3849, 3849, 4095, 4095, 0),
		(drawing, 3850, 3850, 4095, 4095, 0),
		(drawing, 3851, 3851, 4095, 4095, 0),
		(drawing, 3852, 3852, 4095, 4095, 0),
		(drawing, 3853, 3853, 4095, 4095, 0),
		(drawing, 3854, 3854, 4095, 4095, 0),
		(drawing, 3855, 3855, 4095, 4095, 0),
		(drawing, 3856, 3856, 4095, 4095, 0),
		(drawing, 3857, 3857, 4095, 4095, 0),
		(drawing, 3858, 3858, 4095, 4095, 0),
		(drawing, 3859, 3859, 4095, 4095, 0),
		(drawing, 3860, 3860, 4095, 4095, 0),
		(drawing, 3861, 3861, 4095, 4095, 0),
		(drawing, 3862, 3862, 4095, 4095, 0),
		(drawing, 3863, 3863, 4095, 4095, 0),
		(drawing, 3864, 3864, 4095, 4095, 0),
		(drawing, 3865, 3865, 4095, 4095, 0),
		(drawing, 3866, 3866, 4095, 4095, 0),
		(drawing, 3867, 3867, 4095, 4095, 0),
		(drawing, 3868, 3868, 4095, 4095, 0),
		(drawing, 3869, 3869, 4095, 4095, 0),
		(drawing, 3870, 3870, 4095, 4095, 0),
		(drawing, 3871, 3871, 4095, 4095, 0),
		(drawing, 3872, 3872, 4095, 4095, 0),
		(drawing, 3873, 3873, 4095, 4095, 0),
		(drawing, 3874, 3874, 4095, 4095, 0),
		(drawing, 3875, 3875, 4095, 4095, 0),
		(drawing, 3876, 3876, 4095, 4095, 0),
		(drawing, 3877, 3877, 4095, 4095, 0),
		(drawing, 3878, 3878, 4095, 4095, 0),
		(drawing, 3879, 3879, 4095, 4095, 0),
		(drawing, 3880, 3880, 4095, 4095, 0),
		(drawing, 3881, 3881, 4095, 4095, 0),
		(drawing, 3882, 3882, 4095, 4095, 0),
		(drawing, 3883, 3883, 4095, 4095, 0),
		(drawing, 3884, 3884, 4095, 4095, 0),
		(drawing, 3885, 3885, 4095, 4095, 0),
		(drawing, 3886, 3886, 4095, 4095, 0),
		(drawing, 3887, 3887, 4095, 4095, 0),
		(drawing, 3888, 3888, 4095, 4095, 0),
		(drawing, 3889, 3889, 4095, 4095, 0),
		(drawing, 3890, 3890, 4095, 4095, 0),
		(drawing, 3891, 3891, 4095, 4095, 0),
		(drawing, 3892, 3892, 4095, 4095, 0),
		(drawing, 3893, 3893, 4095, 4095, 0),
		(drawing, 3894, 3894, 4095, 4095, 0),
		(drawing, 3895, 3895, 4095, 4095, 0),
		(drawing, 3896, 3896, 4095, 4095, 0),
		(drawing, 3897, 3897, 4095, 4095, 0),
		(drawing, 3898, 3898, 4095, 4095, 0),
		(drawing, 3899, 3899, 4095, 4095, 0),
		(drawing, 3900, 3900, 4095, 4095, 0),
		(drawing, 3901, 3901, 4095, 4095, 0),
		(drawing, 3902, 3902, 4095, 4095, 0),
		(drawing, 3903, 3903, 4095, 4095, 0),
		(drawing, 3904, 3904, 4095, 4095, 0),
		(drawing, 3905, 3905, 4095, 4095, 0),
		(drawing, 3906, 3906, 4095, 4095, 0),
		(drawing, 3907, 3907, 4095, 4095, 0),
		(drawing, 3908, 3908, 4095, 4095, 0),
		(drawing, 3909, 3909, 4095, 4095, 0),
		(drawing, 3910, 3910, 4095, 4095, 0),
		(drawing, 3911, 3911, 4095, 4095, 0),
		(drawing, 3912, 3912, 4095, 4095, 0),
		(drawing, 3913, 3913, 4095, 4095, 0),
		(drawing, 3914, 3914, 4095, 4095, 0),
		(drawing, 3915, 3915, 4095, 4095, 0),
		(drawing, 3916, 3916, 4095, 4095, 0),
		(drawing, 3917, 3917, 4095, 4095, 0),
		(drawing, 3918, 3918, 4095, 4095, 0),
		(drawing, 3919, 3919, 4095, 4095, 0),
		(drawing, 3920, 3920, 4095, 4095, 0),
		(drawing, 3921, 3921, 4095, 4095, 0),
		(drawing, 3922, 3922, 4095, 4095, 0),
		(drawing, 3923, 3923, 4095, 4095, 0),
		(drawing, 3924, 3924, 4095, 4095, 0),
		(drawing, 3925, 3925, 4095, 4095, 0),
		(drawing, 3926, 3926, 4095, 4095, 0),
		(drawing, 3927, 3927, 4095, 4095, 0),
		(drawing, 3928, 3928, 4095, 4095, 0),
		(drawing, 3929, 3929, 4095, 4095, 0),
		(drawing, 3930, 3930, 4095, 4095, 0),
		(drawing, 3931, 3931, 4095, 4095, 0),
		(drawing, 3932, 3932, 4095, 4095, 0),
		(drawing, 3933, 3933, 4095, 4095, 0),
		(drawing, 3934, 3934, 4095, 4095, 0),
		(drawing, 3935, 3935, 4095, 4095, 0),
		(drawing, 3936, 3936, 4095, 4095, 0),
		(drawing, 3937, 3937, 4095, 4095, 0),
		(drawing, 3938, 3938, 4095, 4095, 0),
		(drawing, 3939, 3939, 4095, 4095, 0),
		(drawing, 3940, 3940, 4095, 4095, 0),
		(drawing, 3941, 3941, 4095, 4095, 0),
		(drawing, 3942, 3942, 4095, 4095, 0),
		(drawing, 3943, 3943, 4095, 4095, 0),
		(drawing, 3944, 3944, 4095, 4095, 0),
		(drawing, 3945, 3945, 4095, 4095, 0),
		(drawing, 3946, 3946, 4095, 4095, 0),
		(drawing, 3947, 3947, 4095, 4095, 0),
		(drawing, 3948, 3948, 4095, 4095, 0),
		(drawing, 3949, 3949, 4095, 4095, 0),
		(drawing, 3950, 3950, 4095, 4095, 0),
		(drawing, 3951, 3951, 4095, 4095, 0),
		(drawing, 3952, 3952, 4095, 4095, 0),
		(drawing, 3953, 3953, 4095, 4095, 0),
		(drawing, 3954, 3954, 4095, 4095, 0),
		(drawing, 3955, 3955, 4095, 4095, 0),
		(drawing, 3956, 3956, 4095, 4095, 0),
		(drawing, 3957, 3957, 4095, 4095, 0),
		(drawing, 3958, 3958, 4095, 4095, 0),
		(drawing, 3959, 3959, 4095, 4095, 0),
		(drawing, 3960, 3960, 4095, 4095, 0),
		(drawing, 3961, 3961, 4095, 4095, 0),
		(drawing, 3962, 3962, 4095, 4095, 0),
		(drawing, 3963, 3963, 4095, 4095, 0),
		(drawing, 3964, 3964, 4095, 4095, 0),
		(drawing, 3965, 3965, 4095, 4095, 0),
		(drawing, 3966, 3966, 4095, 4095, 0),
		(drawing, 3967, 3967, 4095, 4095, 0),
		(drawing, 3968, 3968, 4095, 4095, 0),
		(drawing, 3969, 3969, 4095, 4095, 0),
		(drawing, 3970, 3970, 4095, 4095, 0),
		(drawing, 3971, 3971, 4095, 4095, 0),
		(drawing, 3972, 3972, 4095, 4095, 0),
		(drawing, 3973, 3973, 4095, 4095, 0),
		(drawing, 3974, 3974, 4095, 4095, 0),
		(drawing, 3975, 3975, 4095, 4095, 0),
		(drawing, 3976, 3976, 4095, 4095, 0),
		(drawing, 3977, 3977, 4095, 4095, 0),
		(drawing, 3978, 3978, 4095, 4095, 0),
		(drawing, 3979, 3979, 4095, 4095, 0),
		(drawing, 3980, 3980, 4095, 4095, 0),
		(drawing, 3981, 3981, 4095, 4095, 0),
		(drawing, 3982, 3982, 4095, 4095, 0),
		(drawing, 3983, 3983, 4095, 4095, 0),
		(drawing, 3984, 3984, 4095, 4095, 0),
		(drawing, 3985, 3985, 4095, 4095, 0),
		(drawing, 3986, 3986, 4095, 4095, 0),
		(drawing, 3987, 3987, 4095, 4095, 0),
		(drawing, 3988, 3988, 4095, 4095, 0),
		(drawing, 3989, 3989, 4095, 4095, 0),
		(drawing, 3990, 3990, 4095, 4095, 0),
		(drawing, 3991, 3991, 4095, 4095, 0),
		(drawing, 3992, 3992, 4095, 4095, 0),
		(drawing, 3993, 3993, 4095, 4095, 0),
		(drawing, 3994, 3994, 4095, 4095, 0),
		(drawing, 3995, 3995, 4095, 4095, 0),
		(drawing, 3996, 3996, 4095, 4095, 0),
		(drawing, 3997, 3997, 4095, 4095, 0),
		(drawing, 3998, 3998, 4095, 4095, 0),
		(drawing, 3999, 3999, 4095, 4095, 0),
		(drawing, 4000, 4000, 4095, 4095, 0),
		(drawing, 4001, 4001, 4095, 4095, 0),
		(drawing, 4002, 4002, 4095, 4095, 0),
		(drawing, 4003, 4003, 4095, 4095, 0),
		(drawing, 4004, 4004, 4095, 4095, 0),
		(drawing, 4005, 4005, 4095, 4095, 0),
		(drawing, 4006, 4006, 4095, 4095, 0),
		(drawing, 4007, 4007, 4095, 4095, 0),
		(drawing, 4008, 4008, 4095, 4095, 0),
		(drawing, 4009, 4009, 4095, 4095, 0),
		(drawing, 4010, 4010, 4095, 4095, 0),
		(drawing, 4011, 4011, 4095, 4095, 0),
		(drawing, 4012, 4012, 4095, 4095, 0),
		(drawing, 4013, 4013, 4095, 4095, 0),
		(drawing, 4014, 4014, 4095, 4095, 0),
		(drawing, 4015, 4015, 4095, 4095, 0),
		(drawing, 4016, 4016, 4095, 4095, 0),
		(drawing, 4017, 4017, 4095, 4095, 0),
		(drawing, 4018, 4018, 4095, 4095, 0),
		(drawing, 4019, 4019, 4095, 4095, 0),
		(drawing, 4020, 4020, 4095, 4095, 0),
		(drawing, 4021, 4021, 4095, 4095, 0),
		(drawing, 4022, 4022, 4095, 4095, 0),
		(drawing, 4023, 4023, 4095, 4095, 0),
		(drawing, 4024, 4024, 4095, 4095, 0),
		(drawing, 4025, 4025, 4095, 4095, 0),
		(drawing, 4026, 4026, 4095, 4095, 0),
		(drawing, 4027, 4027, 4095, 4095, 0),
		(drawing, 4028, 4028, 4095, 4095, 0),
		(drawing, 4029, 4029, 4095, 4095, 0),
		(drawing, 4030, 4030, 4095, 4095, 0),
		(drawing, 4031, 4031, 4095, 4095, 0),
		(drawing, 4032, 4032, 4095, 4095, 0),
		(drawing, 4033, 4033, 4095, 4095, 0),
		(drawing, 4034, 4034, 4095, 4095, 0),
		(drawing, 4035, 4035, 4095, 4095, 0),
		(drawing, 4036, 4036, 4095, 4095, 0),
		(drawing, 4037, 4037, 4095, 4095, 0),
		(drawing, 4038, 4038, 4095, 4095, 0),
		(drawing, 4039, 4039, 4095, 4095, 0),
		(drawing, 4040, 4040, 4095, 4095, 0),
		(drawing, 4041, 4041, 4095, 4095, 0),
		(drawing, 4042, 4042, 4095, 4095, 0),
		(drawing, 4043, 4043, 4095, 4095, 0),
		(drawing, 4044, 4044, 4095, 4095, 0),
		(drawing, 4045, 4045, 4095, 4095, 0),
		(drawing, 4046, 4046, 4095, 4095, 0),
		(drawing, 4047, 4047, 4095, 4095, 0),
		(drawing, 4048, 4048, 4095, 4095, 0),
		(drawing, 4049, 4049, 4095, 4095, 0),
		(drawing, 4050, 4050, 4095, 4095, 0),
		(drawing, 4051, 4051, 4095, 4095, 0),
		(drawing, 4052, 4052, 4095, 4095, 0),
		(drawing, 4053, 4053, 4095, 4095, 0),
		(drawing, 4054, 4054, 4095, 4095, 0),
		(drawing, 4055, 4055, 4095, 4095, 0),
		(drawing, 4056, 4056, 4095, 4095, 0),
		(drawing, 4057, 4057, 4095, 4095, 0),
		(drawing, 4058, 4058, 4095, 4095, 0),
		(drawing, 4059, 4059, 4095, 4095, 0),
		(drawing, 4060, 4060, 4095, 4095, 0),
		(drawing, 4061, 4061, 4095, 4095, 0),
		(drawing, 4062, 4062, 4095, 4095, 0),
		(drawing, 4063, 4063, 4095, 4095, 0),
		(drawing, 4064, 4064, 4095, 4095, 0),
		(drawing, 4065, 4065, 4095, 4095, 0),
		(drawing, 4066, 4066, 4095, 4095, 0),
		(drawing, 4067, 4067, 4095, 4095, 0),
		(drawing, 4068, 4068, 4095, 4095, 0),
		(drawing, 4069, 4069, 4095, 4095, 0),
		(drawing, 4070, 4070, 4095, 4095, 0),
		(drawing, 4071, 4071, 4095, 4095, 0),
		(drawing, 4072, 4072, 4095, 4095, 0),
		(drawing, 4073, 4073, 4095, 4095, 0),
		(drawing, 4074, 4074, 4095, 4095, 0),
		(drawing, 4075, 4075, 4095, 4095, 0),
		(drawing, 4076, 4076, 4095, 4095, 0),
		(drawing, 4077, 4077, 4095, 4095, 0),
		(drawing, 4078, 4078, 4095, 4095, 0),
		(drawing, 4079, 4079, 4095, 4095, 0),
		(drawing, 4080, 4080, 4095, 4095, 0),
		(drawing, 4081, 4081, 4095, 4095, 0),
		(drawing, 4082, 4082, 4095, 4095, 0),
		(drawing, 4083, 4083, 4095, 4095, 0),
		(drawing, 4084, 4084, 4095, 4095, 0),
		(drawing, 4085, 4085, 4095, 4095, 0),
		(drawing, 4086, 4086, 4095, 4095, 0),
		(drawing, 4087, 4087, 4095, 4095, 0),
		(drawing, 4088, 4088, 4095, 4095, 0),
		(drawing, 4089, 4089, 4095, 4095, 0),
		(drawing, 4090, 4090, 4095, 4095, 0),
		(drawing, 4091, 4091, 4095, 4095, 0),
		(drawing, 4092, 4092, 4095, 4095, 0),
		(drawing, 4093, 4093, 4095, 4095, 0),
		(drawing, 4094, 4094, 4095, 4095, 0),
		(done, 4095, 4095, 4095, 4095, 0)
	);
END PACKAGE ex1_data_pak;
