-- advanced test 9
-- draw line from (35,89) to (3900,800)
-- this is a random test

PACKAGE ex1_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 35, 89, 0),
		(start, 35, 89, 3900, 800, 0),
		(drawing, 35, 89, 3900, 800, 0),
		(drawing, 36, 89, 3900, 800, 0),
		(drawing, 37, 89, 3900, 800, 0),
		(drawing, 38, 90, 3900, 800, 0),
		(drawing, 39, 90, 3900, 800, 0),
		(drawing, 40, 90, 3900, 800, 0),
		(drawing, 41, 90, 3900, 800, 0),
		(drawing, 42, 90, 3900, 800, 0),
		(drawing, 43, 90, 3900, 800, 0),
		(drawing, 44, 91, 3900, 800, 0),
		(drawing, 45, 91, 3900, 800, 0),
		(drawing, 46, 91, 3900, 800, 0),
		(drawing, 47, 91, 3900, 800, 0),
		(drawing, 48, 91, 3900, 800, 0),
		(drawing, 49, 92, 3900, 800, 0),
		(drawing, 50, 92, 3900, 800, 0),
		(drawing, 51, 92, 3900, 800, 0),
		(drawing, 52, 92, 3900, 800, 0),
		(drawing, 53, 92, 3900, 800, 0),
		(drawing, 54, 92, 3900, 800, 0),
		(drawing, 55, 93, 3900, 800, 0),
		(drawing, 56, 93, 3900, 800, 0),
		(drawing, 57, 93, 3900, 800, 0),
		(drawing, 58, 93, 3900, 800, 0),
		(drawing, 59, 93, 3900, 800, 0),
		(drawing, 60, 94, 3900, 800, 0),
		(drawing, 61, 94, 3900, 800, 0),
		(drawing, 62, 94, 3900, 800, 0),
		(drawing, 63, 94, 3900, 800, 0),
		(drawing, 64, 94, 3900, 800, 0),
		(drawing, 65, 95, 3900, 800, 0),
		(drawing, 66, 95, 3900, 800, 0),
		(drawing, 67, 95, 3900, 800, 0),
		(drawing, 68, 95, 3900, 800, 0),
		(drawing, 69, 95, 3900, 800, 0),
		(drawing, 70, 95, 3900, 800, 0),
		(drawing, 71, 96, 3900, 800, 0),
		(drawing, 72, 96, 3900, 800, 0),
		(drawing, 73, 96, 3900, 800, 0),
		(drawing, 74, 96, 3900, 800, 0),
		(drawing, 75, 96, 3900, 800, 0),
		(drawing, 76, 97, 3900, 800, 0),
		(drawing, 77, 97, 3900, 800, 0),
		(drawing, 78, 97, 3900, 800, 0),
		(drawing, 79, 97, 3900, 800, 0),
		(drawing, 80, 97, 3900, 800, 0),
		(drawing, 81, 97, 3900, 800, 0),
		(drawing, 82, 98, 3900, 800, 0),
		(drawing, 83, 98, 3900, 800, 0),
		(drawing, 84, 98, 3900, 800, 0),
		(drawing, 85, 98, 3900, 800, 0),
		(drawing, 86, 98, 3900, 800, 0),
		(drawing, 87, 99, 3900, 800, 0),
		(drawing, 88, 99, 3900, 800, 0),
		(drawing, 89, 99, 3900, 800, 0),
		(drawing, 90, 99, 3900, 800, 0),
		(drawing, 91, 99, 3900, 800, 0),
		(drawing, 92, 99, 3900, 800, 0),
		(drawing, 93, 100, 3900, 800, 0),
		(drawing, 94, 100, 3900, 800, 0),
		(drawing, 95, 100, 3900, 800, 0),
		(drawing, 96, 100, 3900, 800, 0),
		(drawing, 97, 100, 3900, 800, 0),
		(drawing, 98, 101, 3900, 800, 0),
		(drawing, 99, 101, 3900, 800, 0),
		(drawing, 100, 101, 3900, 800, 0),
		(drawing, 101, 101, 3900, 800, 0),
		(drawing, 102, 101, 3900, 800, 0),
		(drawing, 103, 102, 3900, 800, 0),
		(drawing, 104, 102, 3900, 800, 0),
		(drawing, 105, 102, 3900, 800, 0),
		(drawing, 106, 102, 3900, 800, 0),
		(drawing, 107, 102, 3900, 800, 0),
		(drawing, 108, 102, 3900, 800, 0),
		(drawing, 109, 103, 3900, 800, 0),
		(drawing, 110, 103, 3900, 800, 0),
		(drawing, 111, 103, 3900, 800, 0),
		(drawing, 112, 103, 3900, 800, 0),
		(drawing, 113, 103, 3900, 800, 0),
		(drawing, 114, 104, 3900, 800, 0),
		(drawing, 115, 104, 3900, 800, 0),
		(drawing, 116, 104, 3900, 800, 0),
		(drawing, 117, 104, 3900, 800, 0),
		(drawing, 118, 104, 3900, 800, 0),
		(drawing, 119, 104, 3900, 800, 0),
		(drawing, 120, 105, 3900, 800, 0),
		(drawing, 121, 105, 3900, 800, 0),
		(drawing, 122, 105, 3900, 800, 0),
		(drawing, 123, 105, 3900, 800, 0),
		(drawing, 124, 105, 3900, 800, 0),
		(drawing, 125, 106, 3900, 800, 0),
		(drawing, 126, 106, 3900, 800, 0),
		(drawing, 127, 106, 3900, 800, 0),
		(drawing, 128, 106, 3900, 800, 0),
		(drawing, 129, 106, 3900, 800, 0),
		(drawing, 130, 106, 3900, 800, 0),
		(drawing, 131, 107, 3900, 800, 0),
		(drawing, 132, 107, 3900, 800, 0),
		(drawing, 133, 107, 3900, 800, 0),
		(drawing, 134, 107, 3900, 800, 0),
		(drawing, 135, 107, 3900, 800, 0),
		(drawing, 136, 108, 3900, 800, 0),
		(drawing, 137, 108, 3900, 800, 0),
		(drawing, 138, 108, 3900, 800, 0),
		(drawing, 139, 108, 3900, 800, 0),
		(drawing, 140, 108, 3900, 800, 0),
		(drawing, 141, 108, 3900, 800, 0),
		(drawing, 142, 109, 3900, 800, 0),
		(drawing, 143, 109, 3900, 800, 0),
		(drawing, 144, 109, 3900, 800, 0),
		(drawing, 145, 109, 3900, 800, 0),
		(drawing, 146, 109, 3900, 800, 0),
		(drawing, 147, 110, 3900, 800, 0),
		(drawing, 148, 110, 3900, 800, 0),
		(drawing, 149, 110, 3900, 800, 0),
		(drawing, 150, 110, 3900, 800, 0),
		(drawing, 151, 110, 3900, 800, 0),
		(drawing, 152, 111, 3900, 800, 0),
		(drawing, 153, 111, 3900, 800, 0),
		(drawing, 154, 111, 3900, 800, 0),
		(drawing, 155, 111, 3900, 800, 0),
		(drawing, 156, 111, 3900, 800, 0),
		(drawing, 157, 111, 3900, 800, 0),
		(drawing, 158, 112, 3900, 800, 0),
		(drawing, 159, 112, 3900, 800, 0),
		(drawing, 160, 112, 3900, 800, 0),
		(drawing, 161, 112, 3900, 800, 0),
		(drawing, 162, 112, 3900, 800, 0),
		(drawing, 163, 113, 3900, 800, 0),
		(drawing, 164, 113, 3900, 800, 0),
		(drawing, 165, 113, 3900, 800, 0),
		(drawing, 166, 113, 3900, 800, 0),
		(drawing, 167, 113, 3900, 800, 0),
		(drawing, 168, 113, 3900, 800, 0),
		(drawing, 169, 114, 3900, 800, 0),
		(drawing, 170, 114, 3900, 800, 0),
		(drawing, 171, 114, 3900, 800, 0),
		(drawing, 172, 114, 3900, 800, 0),
		(drawing, 173, 114, 3900, 800, 0),
		(drawing, 174, 115, 3900, 800, 0),
		(drawing, 175, 115, 3900, 800, 0),
		(drawing, 176, 115, 3900, 800, 0),
		(drawing, 177, 115, 3900, 800, 0),
		(drawing, 178, 115, 3900, 800, 0),
		(drawing, 179, 115, 3900, 800, 0),
		(drawing, 180, 116, 3900, 800, 0),
		(drawing, 181, 116, 3900, 800, 0),
		(drawing, 182, 116, 3900, 800, 0),
		(drawing, 183, 116, 3900, 800, 0),
		(drawing, 184, 116, 3900, 800, 0),
		(drawing, 185, 117, 3900, 800, 0),
		(drawing, 186, 117, 3900, 800, 0),
		(drawing, 187, 117, 3900, 800, 0),
		(drawing, 188, 117, 3900, 800, 0),
		(drawing, 189, 117, 3900, 800, 0),
		(drawing, 190, 118, 3900, 800, 0),
		(drawing, 191, 118, 3900, 800, 0),
		(drawing, 192, 118, 3900, 800, 0),
		(drawing, 193, 118, 3900, 800, 0),
		(drawing, 194, 118, 3900, 800, 0),
		(drawing, 195, 118, 3900, 800, 0),
		(drawing, 196, 119, 3900, 800, 0),
		(drawing, 197, 119, 3900, 800, 0),
		(drawing, 198, 119, 3900, 800, 0),
		(drawing, 199, 119, 3900, 800, 0),
		(drawing, 200, 119, 3900, 800, 0),
		(drawing, 201, 120, 3900, 800, 0),
		(drawing, 202, 120, 3900, 800, 0),
		(drawing, 203, 120, 3900, 800, 0),
		(drawing, 204, 120, 3900, 800, 0),
		(drawing, 205, 120, 3900, 800, 0),
		(drawing, 206, 120, 3900, 800, 0),
		(drawing, 207, 121, 3900, 800, 0),
		(drawing, 208, 121, 3900, 800, 0),
		(drawing, 209, 121, 3900, 800, 0),
		(drawing, 210, 121, 3900, 800, 0),
		(drawing, 211, 121, 3900, 800, 0),
		(drawing, 212, 122, 3900, 800, 0),
		(drawing, 213, 122, 3900, 800, 0),
		(drawing, 214, 122, 3900, 800, 0),
		(drawing, 215, 122, 3900, 800, 0),
		(drawing, 216, 122, 3900, 800, 0),
		(drawing, 217, 122, 3900, 800, 0),
		(drawing, 218, 123, 3900, 800, 0),
		(drawing, 219, 123, 3900, 800, 0),
		(drawing, 220, 123, 3900, 800, 0),
		(drawing, 221, 123, 3900, 800, 0),
		(drawing, 222, 123, 3900, 800, 0),
		(drawing, 223, 124, 3900, 800, 0),
		(drawing, 224, 124, 3900, 800, 0),
		(drawing, 225, 124, 3900, 800, 0),
		(drawing, 226, 124, 3900, 800, 0),
		(drawing, 227, 124, 3900, 800, 0),
		(drawing, 228, 125, 3900, 800, 0),
		(drawing, 229, 125, 3900, 800, 0),
		(drawing, 230, 125, 3900, 800, 0),
		(drawing, 231, 125, 3900, 800, 0),
		(drawing, 232, 125, 3900, 800, 0),
		(drawing, 233, 125, 3900, 800, 0),
		(drawing, 234, 126, 3900, 800, 0),
		(drawing, 235, 126, 3900, 800, 0),
		(drawing, 236, 126, 3900, 800, 0),
		(drawing, 237, 126, 3900, 800, 0),
		(drawing, 238, 126, 3900, 800, 0),
		(drawing, 239, 127, 3900, 800, 0),
		(drawing, 240, 127, 3900, 800, 0),
		(drawing, 241, 127, 3900, 800, 0),
		(drawing, 242, 127, 3900, 800, 0),
		(drawing, 243, 127, 3900, 800, 0),
		(drawing, 244, 127, 3900, 800, 0),
		(drawing, 245, 128, 3900, 800, 0),
		(drawing, 246, 128, 3900, 800, 0),
		(drawing, 247, 128, 3900, 800, 0),
		(drawing, 248, 128, 3900, 800, 0),
		(drawing, 249, 128, 3900, 800, 0),
		(drawing, 250, 129, 3900, 800, 0),
		(drawing, 251, 129, 3900, 800, 0),
		(drawing, 252, 129, 3900, 800, 0),
		(drawing, 253, 129, 3900, 800, 0),
		(drawing, 254, 129, 3900, 800, 0),
		(drawing, 255, 129, 3900, 800, 0),
		(drawing, 256, 130, 3900, 800, 0),
		(drawing, 257, 130, 3900, 800, 0),
		(drawing, 258, 130, 3900, 800, 0),
		(drawing, 259, 130, 3900, 800, 0),
		(drawing, 260, 130, 3900, 800, 0),
		(drawing, 261, 131, 3900, 800, 0),
		(drawing, 262, 131, 3900, 800, 0),
		(drawing, 263, 131, 3900, 800, 0),
		(drawing, 264, 131, 3900, 800, 0),
		(drawing, 265, 131, 3900, 800, 0),
		(drawing, 266, 131, 3900, 800, 0),
		(drawing, 267, 132, 3900, 800, 0),
		(drawing, 268, 132, 3900, 800, 0),
		(drawing, 269, 132, 3900, 800, 0),
		(drawing, 270, 132, 3900, 800, 0),
		(drawing, 271, 132, 3900, 800, 0),
		(drawing, 272, 133, 3900, 800, 0),
		(drawing, 273, 133, 3900, 800, 0),
		(drawing, 274, 133, 3900, 800, 0),
		(drawing, 275, 133, 3900, 800, 0),
		(drawing, 276, 133, 3900, 800, 0),
		(drawing, 277, 134, 3900, 800, 0),
		(drawing, 278, 134, 3900, 800, 0),
		(drawing, 279, 134, 3900, 800, 0),
		(drawing, 280, 134, 3900, 800, 0),
		(drawing, 281, 134, 3900, 800, 0),
		(drawing, 282, 134, 3900, 800, 0),
		(drawing, 283, 135, 3900, 800, 0),
		(drawing, 284, 135, 3900, 800, 0),
		(drawing, 285, 135, 3900, 800, 0),
		(drawing, 286, 135, 3900, 800, 0),
		(drawing, 287, 135, 3900, 800, 0),
		(drawing, 288, 136, 3900, 800, 0),
		(drawing, 289, 136, 3900, 800, 0),
		(drawing, 290, 136, 3900, 800, 0),
		(drawing, 291, 136, 3900, 800, 0),
		(drawing, 292, 136, 3900, 800, 0),
		(drawing, 293, 136, 3900, 800, 0),
		(drawing, 294, 137, 3900, 800, 0),
		(drawing, 295, 137, 3900, 800, 0),
		(drawing, 296, 137, 3900, 800, 0),
		(drawing, 297, 137, 3900, 800, 0),
		(drawing, 298, 137, 3900, 800, 0),
		(drawing, 299, 138, 3900, 800, 0),
		(drawing, 300, 138, 3900, 800, 0),
		(drawing, 301, 138, 3900, 800, 0),
		(drawing, 302, 138, 3900, 800, 0),
		(drawing, 303, 138, 3900, 800, 0),
		(drawing, 304, 138, 3900, 800, 0),
		(drawing, 305, 139, 3900, 800, 0),
		(drawing, 306, 139, 3900, 800, 0),
		(drawing, 307, 139, 3900, 800, 0),
		(drawing, 308, 139, 3900, 800, 0),
		(drawing, 309, 139, 3900, 800, 0),
		(drawing, 310, 140, 3900, 800, 0),
		(drawing, 311, 140, 3900, 800, 0),
		(drawing, 312, 140, 3900, 800, 0),
		(drawing, 313, 140, 3900, 800, 0),
		(drawing, 314, 140, 3900, 800, 0),
		(drawing, 315, 141, 3900, 800, 0),
		(drawing, 316, 141, 3900, 800, 0),
		(drawing, 317, 141, 3900, 800, 0),
		(drawing, 318, 141, 3900, 800, 0),
		(drawing, 319, 141, 3900, 800, 0),
		(drawing, 320, 141, 3900, 800, 0),
		(drawing, 321, 142, 3900, 800, 0),
		(drawing, 322, 142, 3900, 800, 0),
		(drawing, 323, 142, 3900, 800, 0),
		(drawing, 324, 142, 3900, 800, 0),
		(drawing, 325, 142, 3900, 800, 0),
		(drawing, 326, 143, 3900, 800, 0),
		(drawing, 327, 143, 3900, 800, 0),
		(drawing, 328, 143, 3900, 800, 0),
		(drawing, 329, 143, 3900, 800, 0),
		(drawing, 330, 143, 3900, 800, 0),
		(drawing, 331, 143, 3900, 800, 0),
		(drawing, 332, 144, 3900, 800, 0),
		(drawing, 333, 144, 3900, 800, 0),
		(drawing, 334, 144, 3900, 800, 0),
		(drawing, 335, 144, 3900, 800, 0),
		(drawing, 336, 144, 3900, 800, 0),
		(drawing, 337, 145, 3900, 800, 0),
		(drawing, 338, 145, 3900, 800, 0),
		(drawing, 339, 145, 3900, 800, 0),
		(drawing, 340, 145, 3900, 800, 0),
		(drawing, 341, 145, 3900, 800, 0),
		(drawing, 342, 145, 3900, 800, 0),
		(drawing, 343, 146, 3900, 800, 0),
		(drawing, 344, 146, 3900, 800, 0),
		(drawing, 345, 146, 3900, 800, 0),
		(drawing, 346, 146, 3900, 800, 0),
		(drawing, 347, 146, 3900, 800, 0),
		(drawing, 348, 147, 3900, 800, 0),
		(drawing, 349, 147, 3900, 800, 0),
		(drawing, 350, 147, 3900, 800, 0),
		(drawing, 351, 147, 3900, 800, 0),
		(drawing, 352, 147, 3900, 800, 0),
		(drawing, 353, 147, 3900, 800, 0),
		(drawing, 354, 148, 3900, 800, 0),
		(drawing, 355, 148, 3900, 800, 0),
		(drawing, 356, 148, 3900, 800, 0),
		(drawing, 357, 148, 3900, 800, 0),
		(drawing, 358, 148, 3900, 800, 0),
		(drawing, 359, 149, 3900, 800, 0),
		(drawing, 360, 149, 3900, 800, 0),
		(drawing, 361, 149, 3900, 800, 0),
		(drawing, 362, 149, 3900, 800, 0),
		(drawing, 363, 149, 3900, 800, 0),
		(drawing, 364, 150, 3900, 800, 0),
		(drawing, 365, 150, 3900, 800, 0),
		(drawing, 366, 150, 3900, 800, 0),
		(drawing, 367, 150, 3900, 800, 0),
		(drawing, 368, 150, 3900, 800, 0),
		(drawing, 369, 150, 3900, 800, 0),
		(drawing, 370, 151, 3900, 800, 0),
		(drawing, 371, 151, 3900, 800, 0),
		(drawing, 372, 151, 3900, 800, 0),
		(drawing, 373, 151, 3900, 800, 0),
		(drawing, 374, 151, 3900, 800, 0),
		(drawing, 375, 152, 3900, 800, 0),
		(drawing, 376, 152, 3900, 800, 0),
		(drawing, 377, 152, 3900, 800, 0),
		(drawing, 378, 152, 3900, 800, 0),
		(drawing, 379, 152, 3900, 800, 0),
		(drawing, 380, 152, 3900, 800, 0),
		(drawing, 381, 153, 3900, 800, 0),
		(drawing, 382, 153, 3900, 800, 0),
		(drawing, 383, 153, 3900, 800, 0),
		(drawing, 384, 153, 3900, 800, 0),
		(drawing, 385, 153, 3900, 800, 0),
		(drawing, 386, 154, 3900, 800, 0),
		(drawing, 387, 154, 3900, 800, 0),
		(drawing, 388, 154, 3900, 800, 0),
		(drawing, 389, 154, 3900, 800, 0),
		(drawing, 390, 154, 3900, 800, 0),
		(drawing, 391, 154, 3900, 800, 0),
		(drawing, 392, 155, 3900, 800, 0),
		(drawing, 393, 155, 3900, 800, 0),
		(drawing, 394, 155, 3900, 800, 0),
		(drawing, 395, 155, 3900, 800, 0),
		(drawing, 396, 155, 3900, 800, 0),
		(drawing, 397, 156, 3900, 800, 0),
		(drawing, 398, 156, 3900, 800, 0),
		(drawing, 399, 156, 3900, 800, 0),
		(drawing, 400, 156, 3900, 800, 0),
		(drawing, 401, 156, 3900, 800, 0),
		(drawing, 402, 157, 3900, 800, 0),
		(drawing, 403, 157, 3900, 800, 0),
		(drawing, 404, 157, 3900, 800, 0),
		(drawing, 405, 157, 3900, 800, 0),
		(drawing, 406, 157, 3900, 800, 0),
		(drawing, 407, 157, 3900, 800, 0),
		(drawing, 408, 158, 3900, 800, 0),
		(drawing, 409, 158, 3900, 800, 0),
		(drawing, 410, 158, 3900, 800, 0),
		(drawing, 411, 158, 3900, 800, 0),
		(drawing, 412, 158, 3900, 800, 0),
		(drawing, 413, 159, 3900, 800, 0),
		(drawing, 414, 159, 3900, 800, 0),
		(drawing, 415, 159, 3900, 800, 0),
		(drawing, 416, 159, 3900, 800, 0),
		(drawing, 417, 159, 3900, 800, 0),
		(drawing, 418, 159, 3900, 800, 0),
		(drawing, 419, 160, 3900, 800, 0),
		(drawing, 420, 160, 3900, 800, 0),
		(drawing, 421, 160, 3900, 800, 0),
		(drawing, 422, 160, 3900, 800, 0),
		(drawing, 423, 160, 3900, 800, 0),
		(drawing, 424, 161, 3900, 800, 0),
		(drawing, 425, 161, 3900, 800, 0),
		(drawing, 426, 161, 3900, 800, 0),
		(drawing, 427, 161, 3900, 800, 0),
		(drawing, 428, 161, 3900, 800, 0),
		(drawing, 429, 161, 3900, 800, 0),
		(drawing, 430, 162, 3900, 800, 0),
		(drawing, 431, 162, 3900, 800, 0),
		(drawing, 432, 162, 3900, 800, 0),
		(drawing, 433, 162, 3900, 800, 0),
		(drawing, 434, 162, 3900, 800, 0),
		(drawing, 435, 163, 3900, 800, 0),
		(drawing, 436, 163, 3900, 800, 0),
		(drawing, 437, 163, 3900, 800, 0),
		(drawing, 438, 163, 3900, 800, 0),
		(drawing, 439, 163, 3900, 800, 0),
		(drawing, 440, 164, 3900, 800, 0),
		(drawing, 441, 164, 3900, 800, 0),
		(drawing, 442, 164, 3900, 800, 0),
		(drawing, 443, 164, 3900, 800, 0),
		(drawing, 444, 164, 3900, 800, 0),
		(drawing, 445, 164, 3900, 800, 0),
		(drawing, 446, 165, 3900, 800, 0),
		(drawing, 447, 165, 3900, 800, 0),
		(drawing, 448, 165, 3900, 800, 0),
		(drawing, 449, 165, 3900, 800, 0),
		(drawing, 450, 165, 3900, 800, 0),
		(drawing, 451, 166, 3900, 800, 0),
		(drawing, 452, 166, 3900, 800, 0),
		(drawing, 453, 166, 3900, 800, 0),
		(drawing, 454, 166, 3900, 800, 0),
		(drawing, 455, 166, 3900, 800, 0),
		(drawing, 456, 166, 3900, 800, 0),
		(drawing, 457, 167, 3900, 800, 0),
		(drawing, 458, 167, 3900, 800, 0),
		(drawing, 459, 167, 3900, 800, 0),
		(drawing, 460, 167, 3900, 800, 0),
		(drawing, 461, 167, 3900, 800, 0),
		(drawing, 462, 168, 3900, 800, 0),
		(drawing, 463, 168, 3900, 800, 0),
		(drawing, 464, 168, 3900, 800, 0),
		(drawing, 465, 168, 3900, 800, 0),
		(drawing, 466, 168, 3900, 800, 0),
		(drawing, 467, 168, 3900, 800, 0),
		(drawing, 468, 169, 3900, 800, 0),
		(drawing, 469, 169, 3900, 800, 0),
		(drawing, 470, 169, 3900, 800, 0),
		(drawing, 471, 169, 3900, 800, 0),
		(drawing, 472, 169, 3900, 800, 0),
		(drawing, 473, 170, 3900, 800, 0),
		(drawing, 474, 170, 3900, 800, 0),
		(drawing, 475, 170, 3900, 800, 0),
		(drawing, 476, 170, 3900, 800, 0),
		(drawing, 477, 170, 3900, 800, 0),
		(drawing, 478, 170, 3900, 800, 0),
		(drawing, 479, 171, 3900, 800, 0),
		(drawing, 480, 171, 3900, 800, 0),
		(drawing, 481, 171, 3900, 800, 0),
		(drawing, 482, 171, 3900, 800, 0),
		(drawing, 483, 171, 3900, 800, 0),
		(drawing, 484, 172, 3900, 800, 0),
		(drawing, 485, 172, 3900, 800, 0),
		(drawing, 486, 172, 3900, 800, 0),
		(drawing, 487, 172, 3900, 800, 0),
		(drawing, 488, 172, 3900, 800, 0),
		(drawing, 489, 173, 3900, 800, 0),
		(drawing, 490, 173, 3900, 800, 0),
		(drawing, 491, 173, 3900, 800, 0),
		(drawing, 492, 173, 3900, 800, 0),
		(drawing, 493, 173, 3900, 800, 0),
		(drawing, 494, 173, 3900, 800, 0),
		(drawing, 495, 174, 3900, 800, 0),
		(drawing, 496, 174, 3900, 800, 0),
		(drawing, 497, 174, 3900, 800, 0),
		(drawing, 498, 174, 3900, 800, 0),
		(drawing, 499, 174, 3900, 800, 0),
		(drawing, 500, 175, 3900, 800, 0),
		(drawing, 501, 175, 3900, 800, 0),
		(drawing, 502, 175, 3900, 800, 0),
		(drawing, 503, 175, 3900, 800, 0),
		(drawing, 504, 175, 3900, 800, 0),
		(drawing, 505, 175, 3900, 800, 0),
		(drawing, 506, 176, 3900, 800, 0),
		(drawing, 507, 176, 3900, 800, 0),
		(drawing, 508, 176, 3900, 800, 0),
		(drawing, 509, 176, 3900, 800, 0),
		(drawing, 510, 176, 3900, 800, 0),
		(drawing, 511, 177, 3900, 800, 0),
		(drawing, 512, 177, 3900, 800, 0),
		(drawing, 513, 177, 3900, 800, 0),
		(drawing, 514, 177, 3900, 800, 0),
		(drawing, 515, 177, 3900, 800, 0),
		(drawing, 516, 177, 3900, 800, 0),
		(drawing, 517, 178, 3900, 800, 0),
		(drawing, 518, 178, 3900, 800, 0),
		(drawing, 519, 178, 3900, 800, 0),
		(drawing, 520, 178, 3900, 800, 0),
		(drawing, 521, 178, 3900, 800, 0),
		(drawing, 522, 179, 3900, 800, 0),
		(drawing, 523, 179, 3900, 800, 0),
		(drawing, 524, 179, 3900, 800, 0),
		(drawing, 525, 179, 3900, 800, 0),
		(drawing, 526, 179, 3900, 800, 0),
		(drawing, 527, 180, 3900, 800, 0),
		(drawing, 528, 180, 3900, 800, 0),
		(drawing, 529, 180, 3900, 800, 0),
		(drawing, 530, 180, 3900, 800, 0),
		(drawing, 531, 180, 3900, 800, 0),
		(drawing, 532, 180, 3900, 800, 0),
		(drawing, 533, 181, 3900, 800, 0),
		(drawing, 534, 181, 3900, 800, 0),
		(drawing, 535, 181, 3900, 800, 0),
		(drawing, 536, 181, 3900, 800, 0),
		(drawing, 537, 181, 3900, 800, 0),
		(drawing, 538, 182, 3900, 800, 0),
		(drawing, 539, 182, 3900, 800, 0),
		(drawing, 540, 182, 3900, 800, 0),
		(drawing, 541, 182, 3900, 800, 0),
		(drawing, 542, 182, 3900, 800, 0),
		(drawing, 543, 182, 3900, 800, 0),
		(drawing, 544, 183, 3900, 800, 0),
		(drawing, 545, 183, 3900, 800, 0),
		(drawing, 546, 183, 3900, 800, 0),
		(drawing, 547, 183, 3900, 800, 0),
		(drawing, 548, 183, 3900, 800, 0),
		(drawing, 549, 184, 3900, 800, 0),
		(drawing, 550, 184, 3900, 800, 0),
		(drawing, 551, 184, 3900, 800, 0),
		(drawing, 552, 184, 3900, 800, 0),
		(drawing, 553, 184, 3900, 800, 0),
		(drawing, 554, 184, 3900, 800, 0),
		(drawing, 555, 185, 3900, 800, 0),
		(drawing, 556, 185, 3900, 800, 0),
		(drawing, 557, 185, 3900, 800, 0),
		(drawing, 558, 185, 3900, 800, 0),
		(drawing, 559, 185, 3900, 800, 0),
		(drawing, 560, 186, 3900, 800, 0),
		(drawing, 561, 186, 3900, 800, 0),
		(drawing, 562, 186, 3900, 800, 0),
		(drawing, 563, 186, 3900, 800, 0),
		(drawing, 564, 186, 3900, 800, 0),
		(drawing, 565, 186, 3900, 800, 0),
		(drawing, 566, 187, 3900, 800, 0),
		(drawing, 567, 187, 3900, 800, 0),
		(drawing, 568, 187, 3900, 800, 0),
		(drawing, 569, 187, 3900, 800, 0),
		(drawing, 570, 187, 3900, 800, 0),
		(drawing, 571, 188, 3900, 800, 0),
		(drawing, 572, 188, 3900, 800, 0),
		(drawing, 573, 188, 3900, 800, 0),
		(drawing, 574, 188, 3900, 800, 0),
		(drawing, 575, 188, 3900, 800, 0),
		(drawing, 576, 189, 3900, 800, 0),
		(drawing, 577, 189, 3900, 800, 0),
		(drawing, 578, 189, 3900, 800, 0),
		(drawing, 579, 189, 3900, 800, 0),
		(drawing, 580, 189, 3900, 800, 0),
		(drawing, 581, 189, 3900, 800, 0),
		(drawing, 582, 190, 3900, 800, 0),
		(drawing, 583, 190, 3900, 800, 0),
		(drawing, 584, 190, 3900, 800, 0),
		(drawing, 585, 190, 3900, 800, 0),
		(drawing, 586, 190, 3900, 800, 0),
		(drawing, 587, 191, 3900, 800, 0),
		(drawing, 588, 191, 3900, 800, 0),
		(drawing, 589, 191, 3900, 800, 0),
		(drawing, 590, 191, 3900, 800, 0),
		(drawing, 591, 191, 3900, 800, 0),
		(drawing, 592, 191, 3900, 800, 0),
		(drawing, 593, 192, 3900, 800, 0),
		(drawing, 594, 192, 3900, 800, 0),
		(drawing, 595, 192, 3900, 800, 0),
		(drawing, 596, 192, 3900, 800, 0),
		(drawing, 597, 192, 3900, 800, 0),
		(drawing, 598, 193, 3900, 800, 0),
		(drawing, 599, 193, 3900, 800, 0),
		(drawing, 600, 193, 3900, 800, 0),
		(drawing, 601, 193, 3900, 800, 0),
		(drawing, 602, 193, 3900, 800, 0),
		(drawing, 603, 193, 3900, 800, 0),
		(drawing, 604, 194, 3900, 800, 0),
		(drawing, 605, 194, 3900, 800, 0),
		(drawing, 606, 194, 3900, 800, 0),
		(drawing, 607, 194, 3900, 800, 0),
		(drawing, 608, 194, 3900, 800, 0),
		(drawing, 609, 195, 3900, 800, 0),
		(drawing, 610, 195, 3900, 800, 0),
		(drawing, 611, 195, 3900, 800, 0),
		(drawing, 612, 195, 3900, 800, 0),
		(drawing, 613, 195, 3900, 800, 0),
		(drawing, 614, 196, 3900, 800, 0),
		(drawing, 615, 196, 3900, 800, 0),
		(drawing, 616, 196, 3900, 800, 0),
		(drawing, 617, 196, 3900, 800, 0),
		(drawing, 618, 196, 3900, 800, 0),
		(drawing, 619, 196, 3900, 800, 0),
		(drawing, 620, 197, 3900, 800, 0),
		(drawing, 621, 197, 3900, 800, 0),
		(drawing, 622, 197, 3900, 800, 0),
		(drawing, 623, 197, 3900, 800, 0),
		(drawing, 624, 197, 3900, 800, 0),
		(drawing, 625, 198, 3900, 800, 0),
		(drawing, 626, 198, 3900, 800, 0),
		(drawing, 627, 198, 3900, 800, 0),
		(drawing, 628, 198, 3900, 800, 0),
		(drawing, 629, 198, 3900, 800, 0),
		(drawing, 630, 198, 3900, 800, 0),
		(drawing, 631, 199, 3900, 800, 0),
		(drawing, 632, 199, 3900, 800, 0),
		(drawing, 633, 199, 3900, 800, 0),
		(drawing, 634, 199, 3900, 800, 0),
		(drawing, 635, 199, 3900, 800, 0),
		(drawing, 636, 200, 3900, 800, 0),
		(drawing, 637, 200, 3900, 800, 0),
		(drawing, 638, 200, 3900, 800, 0),
		(drawing, 639, 200, 3900, 800, 0),
		(drawing, 640, 200, 3900, 800, 0),
		(drawing, 641, 200, 3900, 800, 0),
		(drawing, 642, 201, 3900, 800, 0),
		(drawing, 643, 201, 3900, 800, 0),
		(drawing, 644, 201, 3900, 800, 0),
		(drawing, 645, 201, 3900, 800, 0),
		(drawing, 646, 201, 3900, 800, 0),
		(drawing, 647, 202, 3900, 800, 0),
		(drawing, 648, 202, 3900, 800, 0),
		(drawing, 649, 202, 3900, 800, 0),
		(drawing, 650, 202, 3900, 800, 0),
		(drawing, 651, 202, 3900, 800, 0),
		(drawing, 652, 203, 3900, 800, 0),
		(drawing, 653, 203, 3900, 800, 0),
		(drawing, 654, 203, 3900, 800, 0),
		(drawing, 655, 203, 3900, 800, 0),
		(drawing, 656, 203, 3900, 800, 0),
		(drawing, 657, 203, 3900, 800, 0),
		(drawing, 658, 204, 3900, 800, 0),
		(drawing, 659, 204, 3900, 800, 0),
		(drawing, 660, 204, 3900, 800, 0),
		(drawing, 661, 204, 3900, 800, 0),
		(drawing, 662, 204, 3900, 800, 0),
		(drawing, 663, 205, 3900, 800, 0),
		(drawing, 664, 205, 3900, 800, 0),
		(drawing, 665, 205, 3900, 800, 0),
		(drawing, 666, 205, 3900, 800, 0),
		(drawing, 667, 205, 3900, 800, 0),
		(drawing, 668, 205, 3900, 800, 0),
		(drawing, 669, 206, 3900, 800, 0),
		(drawing, 670, 206, 3900, 800, 0),
		(drawing, 671, 206, 3900, 800, 0),
		(drawing, 672, 206, 3900, 800, 0),
		(drawing, 673, 206, 3900, 800, 0),
		(drawing, 674, 207, 3900, 800, 0),
		(drawing, 675, 207, 3900, 800, 0),
		(drawing, 676, 207, 3900, 800, 0),
		(drawing, 677, 207, 3900, 800, 0),
		(drawing, 678, 207, 3900, 800, 0),
		(drawing, 679, 207, 3900, 800, 0),
		(drawing, 680, 208, 3900, 800, 0),
		(drawing, 681, 208, 3900, 800, 0),
		(drawing, 682, 208, 3900, 800, 0),
		(drawing, 683, 208, 3900, 800, 0),
		(drawing, 684, 208, 3900, 800, 0),
		(drawing, 685, 209, 3900, 800, 0),
		(drawing, 686, 209, 3900, 800, 0),
		(drawing, 687, 209, 3900, 800, 0),
		(drawing, 688, 209, 3900, 800, 0),
		(drawing, 689, 209, 3900, 800, 0),
		(drawing, 690, 209, 3900, 800, 0),
		(drawing, 691, 210, 3900, 800, 0),
		(drawing, 692, 210, 3900, 800, 0),
		(drawing, 693, 210, 3900, 800, 0),
		(drawing, 694, 210, 3900, 800, 0),
		(drawing, 695, 210, 3900, 800, 0),
		(drawing, 696, 211, 3900, 800, 0),
		(drawing, 697, 211, 3900, 800, 0),
		(drawing, 698, 211, 3900, 800, 0),
		(drawing, 699, 211, 3900, 800, 0),
		(drawing, 700, 211, 3900, 800, 0),
		(drawing, 701, 212, 3900, 800, 0),
		(drawing, 702, 212, 3900, 800, 0),
		(drawing, 703, 212, 3900, 800, 0),
		(drawing, 704, 212, 3900, 800, 0),
		(drawing, 705, 212, 3900, 800, 0),
		(drawing, 706, 212, 3900, 800, 0),
		(drawing, 707, 213, 3900, 800, 0),
		(drawing, 708, 213, 3900, 800, 0),
		(drawing, 709, 213, 3900, 800, 0),
		(drawing, 710, 213, 3900, 800, 0),
		(drawing, 711, 213, 3900, 800, 0),
		(drawing, 712, 214, 3900, 800, 0),
		(drawing, 713, 214, 3900, 800, 0),
		(drawing, 714, 214, 3900, 800, 0),
		(drawing, 715, 214, 3900, 800, 0),
		(drawing, 716, 214, 3900, 800, 0),
		(drawing, 717, 214, 3900, 800, 0),
		(drawing, 718, 215, 3900, 800, 0),
		(drawing, 719, 215, 3900, 800, 0),
		(drawing, 720, 215, 3900, 800, 0),
		(drawing, 721, 215, 3900, 800, 0),
		(drawing, 722, 215, 3900, 800, 0),
		(drawing, 723, 216, 3900, 800, 0),
		(drawing, 724, 216, 3900, 800, 0),
		(drawing, 725, 216, 3900, 800, 0),
		(drawing, 726, 216, 3900, 800, 0),
		(drawing, 727, 216, 3900, 800, 0),
		(drawing, 728, 216, 3900, 800, 0),
		(drawing, 729, 217, 3900, 800, 0),
		(drawing, 730, 217, 3900, 800, 0),
		(drawing, 731, 217, 3900, 800, 0),
		(drawing, 732, 217, 3900, 800, 0),
		(drawing, 733, 217, 3900, 800, 0),
		(drawing, 734, 218, 3900, 800, 0),
		(drawing, 735, 218, 3900, 800, 0),
		(drawing, 736, 218, 3900, 800, 0),
		(drawing, 737, 218, 3900, 800, 0),
		(drawing, 738, 218, 3900, 800, 0),
		(drawing, 739, 219, 3900, 800, 0),
		(drawing, 740, 219, 3900, 800, 0),
		(drawing, 741, 219, 3900, 800, 0),
		(drawing, 742, 219, 3900, 800, 0),
		(drawing, 743, 219, 3900, 800, 0),
		(drawing, 744, 219, 3900, 800, 0),
		(drawing, 745, 220, 3900, 800, 0),
		(drawing, 746, 220, 3900, 800, 0),
		(drawing, 747, 220, 3900, 800, 0),
		(drawing, 748, 220, 3900, 800, 0),
		(drawing, 749, 220, 3900, 800, 0),
		(drawing, 750, 221, 3900, 800, 0),
		(drawing, 751, 221, 3900, 800, 0),
		(drawing, 752, 221, 3900, 800, 0),
		(drawing, 753, 221, 3900, 800, 0),
		(drawing, 754, 221, 3900, 800, 0),
		(drawing, 755, 221, 3900, 800, 0),
		(drawing, 756, 222, 3900, 800, 0),
		(drawing, 757, 222, 3900, 800, 0),
		(drawing, 758, 222, 3900, 800, 0),
		(drawing, 759, 222, 3900, 800, 0),
		(drawing, 760, 222, 3900, 800, 0),
		(drawing, 761, 223, 3900, 800, 0),
		(drawing, 762, 223, 3900, 800, 0),
		(drawing, 763, 223, 3900, 800, 0),
		(drawing, 764, 223, 3900, 800, 0),
		(drawing, 765, 223, 3900, 800, 0),
		(drawing, 766, 223, 3900, 800, 0),
		(drawing, 767, 224, 3900, 800, 0),
		(drawing, 768, 224, 3900, 800, 0),
		(drawing, 769, 224, 3900, 800, 0),
		(drawing, 770, 224, 3900, 800, 0),
		(drawing, 771, 224, 3900, 800, 0),
		(drawing, 772, 225, 3900, 800, 0),
		(drawing, 773, 225, 3900, 800, 0),
		(drawing, 774, 225, 3900, 800, 0),
		(drawing, 775, 225, 3900, 800, 0),
		(drawing, 776, 225, 3900, 800, 0),
		(drawing, 777, 225, 3900, 800, 0),
		(drawing, 778, 226, 3900, 800, 0),
		(drawing, 779, 226, 3900, 800, 0),
		(drawing, 780, 226, 3900, 800, 0),
		(drawing, 781, 226, 3900, 800, 0),
		(drawing, 782, 226, 3900, 800, 0),
		(drawing, 783, 227, 3900, 800, 0),
		(drawing, 784, 227, 3900, 800, 0),
		(drawing, 785, 227, 3900, 800, 0),
		(drawing, 786, 227, 3900, 800, 0),
		(drawing, 787, 227, 3900, 800, 0),
		(drawing, 788, 228, 3900, 800, 0),
		(drawing, 789, 228, 3900, 800, 0),
		(drawing, 790, 228, 3900, 800, 0),
		(drawing, 791, 228, 3900, 800, 0),
		(drawing, 792, 228, 3900, 800, 0),
		(drawing, 793, 228, 3900, 800, 0),
		(drawing, 794, 229, 3900, 800, 0),
		(drawing, 795, 229, 3900, 800, 0),
		(drawing, 796, 229, 3900, 800, 0),
		(drawing, 797, 229, 3900, 800, 0),
		(drawing, 798, 229, 3900, 800, 0),
		(drawing, 799, 230, 3900, 800, 0),
		(drawing, 800, 230, 3900, 800, 0),
		(drawing, 801, 230, 3900, 800, 0),
		(drawing, 802, 230, 3900, 800, 0),
		(drawing, 803, 230, 3900, 800, 0),
		(drawing, 804, 230, 3900, 800, 0),
		(drawing, 805, 231, 3900, 800, 0),
		(drawing, 806, 231, 3900, 800, 0),
		(drawing, 807, 231, 3900, 800, 0),
		(drawing, 808, 231, 3900, 800, 0),
		(drawing, 809, 231, 3900, 800, 0),
		(drawing, 810, 232, 3900, 800, 0),
		(drawing, 811, 232, 3900, 800, 0),
		(drawing, 812, 232, 3900, 800, 0),
		(drawing, 813, 232, 3900, 800, 0),
		(drawing, 814, 232, 3900, 800, 0),
		(drawing, 815, 232, 3900, 800, 0),
		(drawing, 816, 233, 3900, 800, 0),
		(drawing, 817, 233, 3900, 800, 0),
		(drawing, 818, 233, 3900, 800, 0),
		(drawing, 819, 233, 3900, 800, 0),
		(drawing, 820, 233, 3900, 800, 0),
		(drawing, 821, 234, 3900, 800, 0),
		(drawing, 822, 234, 3900, 800, 0),
		(drawing, 823, 234, 3900, 800, 0),
		(drawing, 824, 234, 3900, 800, 0),
		(drawing, 825, 234, 3900, 800, 0),
		(drawing, 826, 235, 3900, 800, 0),
		(drawing, 827, 235, 3900, 800, 0),
		(drawing, 828, 235, 3900, 800, 0),
		(drawing, 829, 235, 3900, 800, 0),
		(drawing, 830, 235, 3900, 800, 0),
		(drawing, 831, 235, 3900, 800, 0),
		(drawing, 832, 236, 3900, 800, 0),
		(drawing, 833, 236, 3900, 800, 0),
		(drawing, 834, 236, 3900, 800, 0),
		(drawing, 835, 236, 3900, 800, 0),
		(drawing, 836, 236, 3900, 800, 0),
		(drawing, 837, 237, 3900, 800, 0),
		(drawing, 838, 237, 3900, 800, 0),
		(drawing, 839, 237, 3900, 800, 0),
		(drawing, 840, 237, 3900, 800, 0),
		(drawing, 841, 237, 3900, 800, 0),
		(drawing, 842, 237, 3900, 800, 0),
		(drawing, 843, 238, 3900, 800, 0),
		(drawing, 844, 238, 3900, 800, 0),
		(drawing, 845, 238, 3900, 800, 0),
		(drawing, 846, 238, 3900, 800, 0),
		(drawing, 847, 238, 3900, 800, 0),
		(drawing, 848, 239, 3900, 800, 0),
		(drawing, 849, 239, 3900, 800, 0),
		(drawing, 850, 239, 3900, 800, 0),
		(drawing, 851, 239, 3900, 800, 0),
		(drawing, 852, 239, 3900, 800, 0),
		(drawing, 853, 239, 3900, 800, 0),
		(drawing, 854, 240, 3900, 800, 0),
		(drawing, 855, 240, 3900, 800, 0),
		(drawing, 856, 240, 3900, 800, 0),
		(drawing, 857, 240, 3900, 800, 0),
		(drawing, 858, 240, 3900, 800, 0),
		(drawing, 859, 241, 3900, 800, 0),
		(drawing, 860, 241, 3900, 800, 0),
		(drawing, 861, 241, 3900, 800, 0),
		(drawing, 862, 241, 3900, 800, 0),
		(drawing, 863, 241, 3900, 800, 0),
		(drawing, 864, 242, 3900, 800, 0),
		(drawing, 865, 242, 3900, 800, 0),
		(drawing, 866, 242, 3900, 800, 0),
		(drawing, 867, 242, 3900, 800, 0),
		(drawing, 868, 242, 3900, 800, 0),
		(drawing, 869, 242, 3900, 800, 0),
		(drawing, 870, 243, 3900, 800, 0),
		(drawing, 871, 243, 3900, 800, 0),
		(drawing, 872, 243, 3900, 800, 0),
		(drawing, 873, 243, 3900, 800, 0),
		(drawing, 874, 243, 3900, 800, 0),
		(drawing, 875, 244, 3900, 800, 0),
		(drawing, 876, 244, 3900, 800, 0),
		(drawing, 877, 244, 3900, 800, 0),
		(drawing, 878, 244, 3900, 800, 0),
		(drawing, 879, 244, 3900, 800, 0),
		(drawing, 880, 244, 3900, 800, 0),
		(drawing, 881, 245, 3900, 800, 0),
		(drawing, 882, 245, 3900, 800, 0),
		(drawing, 883, 245, 3900, 800, 0),
		(drawing, 884, 245, 3900, 800, 0),
		(drawing, 885, 245, 3900, 800, 0),
		(drawing, 886, 246, 3900, 800, 0),
		(drawing, 887, 246, 3900, 800, 0),
		(drawing, 888, 246, 3900, 800, 0),
		(drawing, 889, 246, 3900, 800, 0),
		(drawing, 890, 246, 3900, 800, 0),
		(drawing, 891, 246, 3900, 800, 0),
		(drawing, 892, 247, 3900, 800, 0),
		(drawing, 893, 247, 3900, 800, 0),
		(drawing, 894, 247, 3900, 800, 0),
		(drawing, 895, 247, 3900, 800, 0),
		(drawing, 896, 247, 3900, 800, 0),
		(drawing, 897, 248, 3900, 800, 0),
		(drawing, 898, 248, 3900, 800, 0),
		(drawing, 899, 248, 3900, 800, 0),
		(drawing, 900, 248, 3900, 800, 0),
		(drawing, 901, 248, 3900, 800, 0),
		(drawing, 902, 248, 3900, 800, 0),
		(drawing, 903, 249, 3900, 800, 0),
		(drawing, 904, 249, 3900, 800, 0),
		(drawing, 905, 249, 3900, 800, 0),
		(drawing, 906, 249, 3900, 800, 0),
		(drawing, 907, 249, 3900, 800, 0),
		(drawing, 908, 250, 3900, 800, 0),
		(drawing, 909, 250, 3900, 800, 0),
		(drawing, 910, 250, 3900, 800, 0),
		(drawing, 911, 250, 3900, 800, 0),
		(drawing, 912, 250, 3900, 800, 0),
		(drawing, 913, 251, 3900, 800, 0),
		(drawing, 914, 251, 3900, 800, 0),
		(drawing, 915, 251, 3900, 800, 0),
		(drawing, 916, 251, 3900, 800, 0),
		(drawing, 917, 251, 3900, 800, 0),
		(drawing, 918, 251, 3900, 800, 0),
		(drawing, 919, 252, 3900, 800, 0),
		(drawing, 920, 252, 3900, 800, 0),
		(drawing, 921, 252, 3900, 800, 0),
		(drawing, 922, 252, 3900, 800, 0),
		(drawing, 923, 252, 3900, 800, 0),
		(drawing, 924, 253, 3900, 800, 0),
		(drawing, 925, 253, 3900, 800, 0),
		(drawing, 926, 253, 3900, 800, 0),
		(drawing, 927, 253, 3900, 800, 0),
		(drawing, 928, 253, 3900, 800, 0),
		(drawing, 929, 253, 3900, 800, 0),
		(drawing, 930, 254, 3900, 800, 0),
		(drawing, 931, 254, 3900, 800, 0),
		(drawing, 932, 254, 3900, 800, 0),
		(drawing, 933, 254, 3900, 800, 0),
		(drawing, 934, 254, 3900, 800, 0),
		(drawing, 935, 255, 3900, 800, 0),
		(drawing, 936, 255, 3900, 800, 0),
		(drawing, 937, 255, 3900, 800, 0),
		(drawing, 938, 255, 3900, 800, 0),
		(drawing, 939, 255, 3900, 800, 0),
		(drawing, 940, 255, 3900, 800, 0),
		(drawing, 941, 256, 3900, 800, 0),
		(drawing, 942, 256, 3900, 800, 0),
		(drawing, 943, 256, 3900, 800, 0),
		(drawing, 944, 256, 3900, 800, 0),
		(drawing, 945, 256, 3900, 800, 0),
		(drawing, 946, 257, 3900, 800, 0),
		(drawing, 947, 257, 3900, 800, 0),
		(drawing, 948, 257, 3900, 800, 0),
		(drawing, 949, 257, 3900, 800, 0),
		(drawing, 950, 257, 3900, 800, 0),
		(drawing, 951, 258, 3900, 800, 0),
		(drawing, 952, 258, 3900, 800, 0),
		(drawing, 953, 258, 3900, 800, 0),
		(drawing, 954, 258, 3900, 800, 0),
		(drawing, 955, 258, 3900, 800, 0),
		(drawing, 956, 258, 3900, 800, 0),
		(drawing, 957, 259, 3900, 800, 0),
		(drawing, 958, 259, 3900, 800, 0),
		(drawing, 959, 259, 3900, 800, 0),
		(drawing, 960, 259, 3900, 800, 0),
		(drawing, 961, 259, 3900, 800, 0),
		(drawing, 962, 260, 3900, 800, 0),
		(drawing, 963, 260, 3900, 800, 0),
		(drawing, 964, 260, 3900, 800, 0),
		(drawing, 965, 260, 3900, 800, 0),
		(drawing, 966, 260, 3900, 800, 0),
		(drawing, 967, 260, 3900, 800, 0),
		(drawing, 968, 261, 3900, 800, 0),
		(drawing, 969, 261, 3900, 800, 0),
		(drawing, 970, 261, 3900, 800, 0),
		(drawing, 971, 261, 3900, 800, 0),
		(drawing, 972, 261, 3900, 800, 0),
		(drawing, 973, 262, 3900, 800, 0),
		(drawing, 974, 262, 3900, 800, 0),
		(drawing, 975, 262, 3900, 800, 0),
		(drawing, 976, 262, 3900, 800, 0),
		(drawing, 977, 262, 3900, 800, 0),
		(drawing, 978, 262, 3900, 800, 0),
		(drawing, 979, 263, 3900, 800, 0),
		(drawing, 980, 263, 3900, 800, 0),
		(drawing, 981, 263, 3900, 800, 0),
		(drawing, 982, 263, 3900, 800, 0),
		(drawing, 983, 263, 3900, 800, 0),
		(drawing, 984, 264, 3900, 800, 0),
		(drawing, 985, 264, 3900, 800, 0),
		(drawing, 986, 264, 3900, 800, 0),
		(drawing, 987, 264, 3900, 800, 0),
		(drawing, 988, 264, 3900, 800, 0),
		(drawing, 989, 264, 3900, 800, 0),
		(drawing, 990, 265, 3900, 800, 0),
		(drawing, 991, 265, 3900, 800, 0),
		(drawing, 992, 265, 3900, 800, 0),
		(drawing, 993, 265, 3900, 800, 0),
		(drawing, 994, 265, 3900, 800, 0),
		(drawing, 995, 266, 3900, 800, 0),
		(drawing, 996, 266, 3900, 800, 0),
		(drawing, 997, 266, 3900, 800, 0),
		(drawing, 998, 266, 3900, 800, 0),
		(drawing, 999, 266, 3900, 800, 0),
		(drawing, 1000, 267, 3900, 800, 0),
		(drawing, 1001, 267, 3900, 800, 0),
		(drawing, 1002, 267, 3900, 800, 0),
		(drawing, 1003, 267, 3900, 800, 0),
		(drawing, 1004, 267, 3900, 800, 0),
		(drawing, 1005, 267, 3900, 800, 0),
		(drawing, 1006, 268, 3900, 800, 0),
		(drawing, 1007, 268, 3900, 800, 0),
		(drawing, 1008, 268, 3900, 800, 0),
		(drawing, 1009, 268, 3900, 800, 0),
		(drawing, 1010, 268, 3900, 800, 0),
		(drawing, 1011, 269, 3900, 800, 0),
		(drawing, 1012, 269, 3900, 800, 0),
		(drawing, 1013, 269, 3900, 800, 0),
		(drawing, 1014, 269, 3900, 800, 0),
		(drawing, 1015, 269, 3900, 800, 0),
		(drawing, 1016, 269, 3900, 800, 0),
		(drawing, 1017, 270, 3900, 800, 0),
		(drawing, 1018, 270, 3900, 800, 0),
		(drawing, 1019, 270, 3900, 800, 0),
		(drawing, 1020, 270, 3900, 800, 0),
		(drawing, 1021, 270, 3900, 800, 0),
		(drawing, 1022, 271, 3900, 800, 0),
		(drawing, 1023, 271, 3900, 800, 0),
		(drawing, 1024, 271, 3900, 800, 0),
		(drawing, 1025, 271, 3900, 800, 0),
		(drawing, 1026, 271, 3900, 800, 0),
		(drawing, 1027, 271, 3900, 800, 0),
		(drawing, 1028, 272, 3900, 800, 0),
		(drawing, 1029, 272, 3900, 800, 0),
		(drawing, 1030, 272, 3900, 800, 0),
		(drawing, 1031, 272, 3900, 800, 0),
		(drawing, 1032, 272, 3900, 800, 0),
		(drawing, 1033, 273, 3900, 800, 0),
		(drawing, 1034, 273, 3900, 800, 0),
		(drawing, 1035, 273, 3900, 800, 0),
		(drawing, 1036, 273, 3900, 800, 0),
		(drawing, 1037, 273, 3900, 800, 0),
		(drawing, 1038, 274, 3900, 800, 0),
		(drawing, 1039, 274, 3900, 800, 0),
		(drawing, 1040, 274, 3900, 800, 0),
		(drawing, 1041, 274, 3900, 800, 0),
		(drawing, 1042, 274, 3900, 800, 0),
		(drawing, 1043, 274, 3900, 800, 0),
		(drawing, 1044, 275, 3900, 800, 0),
		(drawing, 1045, 275, 3900, 800, 0),
		(drawing, 1046, 275, 3900, 800, 0),
		(drawing, 1047, 275, 3900, 800, 0),
		(drawing, 1048, 275, 3900, 800, 0),
		(drawing, 1049, 276, 3900, 800, 0),
		(drawing, 1050, 276, 3900, 800, 0),
		(drawing, 1051, 276, 3900, 800, 0),
		(drawing, 1052, 276, 3900, 800, 0),
		(drawing, 1053, 276, 3900, 800, 0),
		(drawing, 1054, 276, 3900, 800, 0),
		(drawing, 1055, 277, 3900, 800, 0),
		(drawing, 1056, 277, 3900, 800, 0),
		(drawing, 1057, 277, 3900, 800, 0),
		(drawing, 1058, 277, 3900, 800, 0),
		(drawing, 1059, 277, 3900, 800, 0),
		(drawing, 1060, 278, 3900, 800, 0),
		(drawing, 1061, 278, 3900, 800, 0),
		(drawing, 1062, 278, 3900, 800, 0),
		(drawing, 1063, 278, 3900, 800, 0),
		(drawing, 1064, 278, 3900, 800, 0),
		(drawing, 1065, 278, 3900, 800, 0),
		(drawing, 1066, 279, 3900, 800, 0),
		(drawing, 1067, 279, 3900, 800, 0),
		(drawing, 1068, 279, 3900, 800, 0),
		(drawing, 1069, 279, 3900, 800, 0),
		(drawing, 1070, 279, 3900, 800, 0),
		(drawing, 1071, 280, 3900, 800, 0),
		(drawing, 1072, 280, 3900, 800, 0),
		(drawing, 1073, 280, 3900, 800, 0),
		(drawing, 1074, 280, 3900, 800, 0),
		(drawing, 1075, 280, 3900, 800, 0),
		(drawing, 1076, 281, 3900, 800, 0),
		(drawing, 1077, 281, 3900, 800, 0),
		(drawing, 1078, 281, 3900, 800, 0),
		(drawing, 1079, 281, 3900, 800, 0),
		(drawing, 1080, 281, 3900, 800, 0),
		(drawing, 1081, 281, 3900, 800, 0),
		(drawing, 1082, 282, 3900, 800, 0),
		(drawing, 1083, 282, 3900, 800, 0),
		(drawing, 1084, 282, 3900, 800, 0),
		(drawing, 1085, 282, 3900, 800, 0),
		(drawing, 1086, 282, 3900, 800, 0),
		(drawing, 1087, 283, 3900, 800, 0),
		(drawing, 1088, 283, 3900, 800, 0),
		(drawing, 1089, 283, 3900, 800, 0),
		(drawing, 1090, 283, 3900, 800, 0),
		(drawing, 1091, 283, 3900, 800, 0),
		(drawing, 1092, 283, 3900, 800, 0),
		(drawing, 1093, 284, 3900, 800, 0),
		(drawing, 1094, 284, 3900, 800, 0),
		(drawing, 1095, 284, 3900, 800, 0),
		(drawing, 1096, 284, 3900, 800, 0),
		(drawing, 1097, 284, 3900, 800, 0),
		(drawing, 1098, 285, 3900, 800, 0),
		(drawing, 1099, 285, 3900, 800, 0),
		(drawing, 1100, 285, 3900, 800, 0),
		(drawing, 1101, 285, 3900, 800, 0),
		(drawing, 1102, 285, 3900, 800, 0),
		(drawing, 1103, 285, 3900, 800, 0),
		(drawing, 1104, 286, 3900, 800, 0),
		(drawing, 1105, 286, 3900, 800, 0),
		(drawing, 1106, 286, 3900, 800, 0),
		(drawing, 1107, 286, 3900, 800, 0),
		(drawing, 1108, 286, 3900, 800, 0),
		(drawing, 1109, 287, 3900, 800, 0),
		(drawing, 1110, 287, 3900, 800, 0),
		(drawing, 1111, 287, 3900, 800, 0),
		(drawing, 1112, 287, 3900, 800, 0),
		(drawing, 1113, 287, 3900, 800, 0),
		(drawing, 1114, 287, 3900, 800, 0),
		(drawing, 1115, 288, 3900, 800, 0),
		(drawing, 1116, 288, 3900, 800, 0),
		(drawing, 1117, 288, 3900, 800, 0),
		(drawing, 1118, 288, 3900, 800, 0),
		(drawing, 1119, 288, 3900, 800, 0),
		(drawing, 1120, 289, 3900, 800, 0),
		(drawing, 1121, 289, 3900, 800, 0),
		(drawing, 1122, 289, 3900, 800, 0),
		(drawing, 1123, 289, 3900, 800, 0),
		(drawing, 1124, 289, 3900, 800, 0),
		(drawing, 1125, 290, 3900, 800, 0),
		(drawing, 1126, 290, 3900, 800, 0),
		(drawing, 1127, 290, 3900, 800, 0),
		(drawing, 1128, 290, 3900, 800, 0),
		(drawing, 1129, 290, 3900, 800, 0),
		(drawing, 1130, 290, 3900, 800, 0),
		(drawing, 1131, 291, 3900, 800, 0),
		(drawing, 1132, 291, 3900, 800, 0),
		(drawing, 1133, 291, 3900, 800, 0),
		(drawing, 1134, 291, 3900, 800, 0),
		(drawing, 1135, 291, 3900, 800, 0),
		(drawing, 1136, 292, 3900, 800, 0),
		(drawing, 1137, 292, 3900, 800, 0),
		(drawing, 1138, 292, 3900, 800, 0),
		(drawing, 1139, 292, 3900, 800, 0),
		(drawing, 1140, 292, 3900, 800, 0),
		(drawing, 1141, 292, 3900, 800, 0),
		(drawing, 1142, 293, 3900, 800, 0),
		(drawing, 1143, 293, 3900, 800, 0),
		(drawing, 1144, 293, 3900, 800, 0),
		(drawing, 1145, 293, 3900, 800, 0),
		(drawing, 1146, 293, 3900, 800, 0),
		(drawing, 1147, 294, 3900, 800, 0),
		(drawing, 1148, 294, 3900, 800, 0),
		(drawing, 1149, 294, 3900, 800, 0),
		(drawing, 1150, 294, 3900, 800, 0),
		(drawing, 1151, 294, 3900, 800, 0),
		(drawing, 1152, 294, 3900, 800, 0),
		(drawing, 1153, 295, 3900, 800, 0),
		(drawing, 1154, 295, 3900, 800, 0),
		(drawing, 1155, 295, 3900, 800, 0),
		(drawing, 1156, 295, 3900, 800, 0),
		(drawing, 1157, 295, 3900, 800, 0),
		(drawing, 1158, 296, 3900, 800, 0),
		(drawing, 1159, 296, 3900, 800, 0),
		(drawing, 1160, 296, 3900, 800, 0),
		(drawing, 1161, 296, 3900, 800, 0),
		(drawing, 1162, 296, 3900, 800, 0),
		(drawing, 1163, 297, 3900, 800, 0),
		(drawing, 1164, 297, 3900, 800, 0),
		(drawing, 1165, 297, 3900, 800, 0),
		(drawing, 1166, 297, 3900, 800, 0),
		(drawing, 1167, 297, 3900, 800, 0),
		(drawing, 1168, 297, 3900, 800, 0),
		(drawing, 1169, 298, 3900, 800, 0),
		(drawing, 1170, 298, 3900, 800, 0),
		(drawing, 1171, 298, 3900, 800, 0),
		(drawing, 1172, 298, 3900, 800, 0),
		(drawing, 1173, 298, 3900, 800, 0),
		(drawing, 1174, 299, 3900, 800, 0),
		(drawing, 1175, 299, 3900, 800, 0),
		(drawing, 1176, 299, 3900, 800, 0),
		(drawing, 1177, 299, 3900, 800, 0),
		(drawing, 1178, 299, 3900, 800, 0),
		(drawing, 1179, 299, 3900, 800, 0),
		(drawing, 1180, 300, 3900, 800, 0),
		(drawing, 1181, 300, 3900, 800, 0),
		(drawing, 1182, 300, 3900, 800, 0),
		(drawing, 1183, 300, 3900, 800, 0),
		(drawing, 1184, 300, 3900, 800, 0),
		(drawing, 1185, 301, 3900, 800, 0),
		(drawing, 1186, 301, 3900, 800, 0),
		(drawing, 1187, 301, 3900, 800, 0),
		(drawing, 1188, 301, 3900, 800, 0),
		(drawing, 1189, 301, 3900, 800, 0),
		(drawing, 1190, 301, 3900, 800, 0),
		(drawing, 1191, 302, 3900, 800, 0),
		(drawing, 1192, 302, 3900, 800, 0),
		(drawing, 1193, 302, 3900, 800, 0),
		(drawing, 1194, 302, 3900, 800, 0),
		(drawing, 1195, 302, 3900, 800, 0),
		(drawing, 1196, 303, 3900, 800, 0),
		(drawing, 1197, 303, 3900, 800, 0),
		(drawing, 1198, 303, 3900, 800, 0),
		(drawing, 1199, 303, 3900, 800, 0),
		(drawing, 1200, 303, 3900, 800, 0),
		(drawing, 1201, 303, 3900, 800, 0),
		(drawing, 1202, 304, 3900, 800, 0),
		(drawing, 1203, 304, 3900, 800, 0),
		(drawing, 1204, 304, 3900, 800, 0),
		(drawing, 1205, 304, 3900, 800, 0),
		(drawing, 1206, 304, 3900, 800, 0),
		(drawing, 1207, 305, 3900, 800, 0),
		(drawing, 1208, 305, 3900, 800, 0),
		(drawing, 1209, 305, 3900, 800, 0),
		(drawing, 1210, 305, 3900, 800, 0),
		(drawing, 1211, 305, 3900, 800, 0),
		(drawing, 1212, 306, 3900, 800, 0),
		(drawing, 1213, 306, 3900, 800, 0),
		(drawing, 1214, 306, 3900, 800, 0),
		(drawing, 1215, 306, 3900, 800, 0),
		(drawing, 1216, 306, 3900, 800, 0),
		(drawing, 1217, 306, 3900, 800, 0),
		(drawing, 1218, 307, 3900, 800, 0),
		(drawing, 1219, 307, 3900, 800, 0),
		(drawing, 1220, 307, 3900, 800, 0),
		(drawing, 1221, 307, 3900, 800, 0),
		(drawing, 1222, 307, 3900, 800, 0),
		(drawing, 1223, 308, 3900, 800, 0),
		(drawing, 1224, 308, 3900, 800, 0),
		(drawing, 1225, 308, 3900, 800, 0),
		(drawing, 1226, 308, 3900, 800, 0),
		(drawing, 1227, 308, 3900, 800, 0),
		(drawing, 1228, 308, 3900, 800, 0),
		(drawing, 1229, 309, 3900, 800, 0),
		(drawing, 1230, 309, 3900, 800, 0),
		(drawing, 1231, 309, 3900, 800, 0),
		(drawing, 1232, 309, 3900, 800, 0),
		(drawing, 1233, 309, 3900, 800, 0),
		(drawing, 1234, 310, 3900, 800, 0),
		(drawing, 1235, 310, 3900, 800, 0),
		(drawing, 1236, 310, 3900, 800, 0),
		(drawing, 1237, 310, 3900, 800, 0),
		(drawing, 1238, 310, 3900, 800, 0),
		(drawing, 1239, 310, 3900, 800, 0),
		(drawing, 1240, 311, 3900, 800, 0),
		(drawing, 1241, 311, 3900, 800, 0),
		(drawing, 1242, 311, 3900, 800, 0),
		(drawing, 1243, 311, 3900, 800, 0),
		(drawing, 1244, 311, 3900, 800, 0),
		(drawing, 1245, 312, 3900, 800, 0),
		(drawing, 1246, 312, 3900, 800, 0),
		(drawing, 1247, 312, 3900, 800, 0),
		(drawing, 1248, 312, 3900, 800, 0),
		(drawing, 1249, 312, 3900, 800, 0),
		(drawing, 1250, 313, 3900, 800, 0),
		(drawing, 1251, 313, 3900, 800, 0),
		(drawing, 1252, 313, 3900, 800, 0),
		(drawing, 1253, 313, 3900, 800, 0),
		(drawing, 1254, 313, 3900, 800, 0),
		(drawing, 1255, 313, 3900, 800, 0),
		(drawing, 1256, 314, 3900, 800, 0),
		(drawing, 1257, 314, 3900, 800, 0),
		(drawing, 1258, 314, 3900, 800, 0),
		(drawing, 1259, 314, 3900, 800, 0),
		(drawing, 1260, 314, 3900, 800, 0),
		(drawing, 1261, 315, 3900, 800, 0),
		(drawing, 1262, 315, 3900, 800, 0),
		(drawing, 1263, 315, 3900, 800, 0),
		(drawing, 1264, 315, 3900, 800, 0),
		(drawing, 1265, 315, 3900, 800, 0),
		(drawing, 1266, 315, 3900, 800, 0),
		(drawing, 1267, 316, 3900, 800, 0),
		(drawing, 1268, 316, 3900, 800, 0),
		(drawing, 1269, 316, 3900, 800, 0),
		(drawing, 1270, 316, 3900, 800, 0),
		(drawing, 1271, 316, 3900, 800, 0),
		(drawing, 1272, 317, 3900, 800, 0),
		(drawing, 1273, 317, 3900, 800, 0),
		(drawing, 1274, 317, 3900, 800, 0),
		(drawing, 1275, 317, 3900, 800, 0),
		(drawing, 1276, 317, 3900, 800, 0),
		(drawing, 1277, 317, 3900, 800, 0),
		(drawing, 1278, 318, 3900, 800, 0),
		(drawing, 1279, 318, 3900, 800, 0),
		(drawing, 1280, 318, 3900, 800, 0),
		(drawing, 1281, 318, 3900, 800, 0),
		(drawing, 1282, 318, 3900, 800, 0),
		(drawing, 1283, 319, 3900, 800, 0),
		(drawing, 1284, 319, 3900, 800, 0),
		(drawing, 1285, 319, 3900, 800, 0),
		(drawing, 1286, 319, 3900, 800, 0),
		(drawing, 1287, 319, 3900, 800, 0),
		(drawing, 1288, 320, 3900, 800, 0),
		(drawing, 1289, 320, 3900, 800, 0),
		(drawing, 1290, 320, 3900, 800, 0),
		(drawing, 1291, 320, 3900, 800, 0),
		(drawing, 1292, 320, 3900, 800, 0),
		(drawing, 1293, 320, 3900, 800, 0),
		(drawing, 1294, 321, 3900, 800, 0),
		(drawing, 1295, 321, 3900, 800, 0),
		(drawing, 1296, 321, 3900, 800, 0),
		(drawing, 1297, 321, 3900, 800, 0),
		(drawing, 1298, 321, 3900, 800, 0),
		(drawing, 1299, 322, 3900, 800, 0),
		(drawing, 1300, 322, 3900, 800, 0),
		(drawing, 1301, 322, 3900, 800, 0),
		(drawing, 1302, 322, 3900, 800, 0),
		(drawing, 1303, 322, 3900, 800, 0),
		(drawing, 1304, 322, 3900, 800, 0),
		(drawing, 1305, 323, 3900, 800, 0),
		(drawing, 1306, 323, 3900, 800, 0),
		(drawing, 1307, 323, 3900, 800, 0),
		(drawing, 1308, 323, 3900, 800, 0),
		(drawing, 1309, 323, 3900, 800, 0),
		(drawing, 1310, 324, 3900, 800, 0),
		(drawing, 1311, 324, 3900, 800, 0),
		(drawing, 1312, 324, 3900, 800, 0),
		(drawing, 1313, 324, 3900, 800, 0),
		(drawing, 1314, 324, 3900, 800, 0),
		(drawing, 1315, 324, 3900, 800, 0),
		(drawing, 1316, 325, 3900, 800, 0),
		(drawing, 1317, 325, 3900, 800, 0),
		(drawing, 1318, 325, 3900, 800, 0),
		(drawing, 1319, 325, 3900, 800, 0),
		(drawing, 1320, 325, 3900, 800, 0),
		(drawing, 1321, 326, 3900, 800, 0),
		(drawing, 1322, 326, 3900, 800, 0),
		(drawing, 1323, 326, 3900, 800, 0),
		(drawing, 1324, 326, 3900, 800, 0),
		(drawing, 1325, 326, 3900, 800, 0),
		(drawing, 1326, 326, 3900, 800, 0),
		(drawing, 1327, 327, 3900, 800, 0),
		(drawing, 1328, 327, 3900, 800, 0),
		(drawing, 1329, 327, 3900, 800, 0),
		(drawing, 1330, 327, 3900, 800, 0),
		(drawing, 1331, 327, 3900, 800, 0),
		(drawing, 1332, 328, 3900, 800, 0),
		(drawing, 1333, 328, 3900, 800, 0),
		(drawing, 1334, 328, 3900, 800, 0),
		(drawing, 1335, 328, 3900, 800, 0),
		(drawing, 1336, 328, 3900, 800, 0),
		(drawing, 1337, 329, 3900, 800, 0),
		(drawing, 1338, 329, 3900, 800, 0),
		(drawing, 1339, 329, 3900, 800, 0),
		(drawing, 1340, 329, 3900, 800, 0),
		(drawing, 1341, 329, 3900, 800, 0),
		(drawing, 1342, 329, 3900, 800, 0),
		(drawing, 1343, 330, 3900, 800, 0),
		(drawing, 1344, 330, 3900, 800, 0),
		(drawing, 1345, 330, 3900, 800, 0),
		(drawing, 1346, 330, 3900, 800, 0),
		(drawing, 1347, 330, 3900, 800, 0),
		(drawing, 1348, 331, 3900, 800, 0),
		(drawing, 1349, 331, 3900, 800, 0),
		(drawing, 1350, 331, 3900, 800, 0),
		(drawing, 1351, 331, 3900, 800, 0),
		(drawing, 1352, 331, 3900, 800, 0),
		(drawing, 1353, 331, 3900, 800, 0),
		(drawing, 1354, 332, 3900, 800, 0),
		(drawing, 1355, 332, 3900, 800, 0),
		(drawing, 1356, 332, 3900, 800, 0),
		(drawing, 1357, 332, 3900, 800, 0),
		(drawing, 1358, 332, 3900, 800, 0),
		(drawing, 1359, 333, 3900, 800, 0),
		(drawing, 1360, 333, 3900, 800, 0),
		(drawing, 1361, 333, 3900, 800, 0),
		(drawing, 1362, 333, 3900, 800, 0),
		(drawing, 1363, 333, 3900, 800, 0),
		(drawing, 1364, 333, 3900, 800, 0),
		(drawing, 1365, 334, 3900, 800, 0),
		(drawing, 1366, 334, 3900, 800, 0),
		(drawing, 1367, 334, 3900, 800, 0),
		(drawing, 1368, 334, 3900, 800, 0),
		(drawing, 1369, 334, 3900, 800, 0),
		(drawing, 1370, 335, 3900, 800, 0),
		(drawing, 1371, 335, 3900, 800, 0),
		(drawing, 1372, 335, 3900, 800, 0),
		(drawing, 1373, 335, 3900, 800, 0),
		(drawing, 1374, 335, 3900, 800, 0),
		(drawing, 1375, 336, 3900, 800, 0),
		(drawing, 1376, 336, 3900, 800, 0),
		(drawing, 1377, 336, 3900, 800, 0),
		(drawing, 1378, 336, 3900, 800, 0),
		(drawing, 1379, 336, 3900, 800, 0),
		(drawing, 1380, 336, 3900, 800, 0),
		(drawing, 1381, 337, 3900, 800, 0),
		(drawing, 1382, 337, 3900, 800, 0),
		(drawing, 1383, 337, 3900, 800, 0),
		(drawing, 1384, 337, 3900, 800, 0),
		(drawing, 1385, 337, 3900, 800, 0),
		(drawing, 1386, 338, 3900, 800, 0),
		(drawing, 1387, 338, 3900, 800, 0),
		(drawing, 1388, 338, 3900, 800, 0),
		(drawing, 1389, 338, 3900, 800, 0),
		(drawing, 1390, 338, 3900, 800, 0),
		(drawing, 1391, 338, 3900, 800, 0),
		(drawing, 1392, 339, 3900, 800, 0),
		(drawing, 1393, 339, 3900, 800, 0),
		(drawing, 1394, 339, 3900, 800, 0),
		(drawing, 1395, 339, 3900, 800, 0),
		(drawing, 1396, 339, 3900, 800, 0),
		(drawing, 1397, 340, 3900, 800, 0),
		(drawing, 1398, 340, 3900, 800, 0),
		(drawing, 1399, 340, 3900, 800, 0),
		(drawing, 1400, 340, 3900, 800, 0),
		(drawing, 1401, 340, 3900, 800, 0),
		(drawing, 1402, 340, 3900, 800, 0),
		(drawing, 1403, 341, 3900, 800, 0),
		(drawing, 1404, 341, 3900, 800, 0),
		(drawing, 1405, 341, 3900, 800, 0),
		(drawing, 1406, 341, 3900, 800, 0),
		(drawing, 1407, 341, 3900, 800, 0),
		(drawing, 1408, 342, 3900, 800, 0),
		(drawing, 1409, 342, 3900, 800, 0),
		(drawing, 1410, 342, 3900, 800, 0),
		(drawing, 1411, 342, 3900, 800, 0),
		(drawing, 1412, 342, 3900, 800, 0),
		(drawing, 1413, 342, 3900, 800, 0),
		(drawing, 1414, 343, 3900, 800, 0),
		(drawing, 1415, 343, 3900, 800, 0),
		(drawing, 1416, 343, 3900, 800, 0),
		(drawing, 1417, 343, 3900, 800, 0),
		(drawing, 1418, 343, 3900, 800, 0),
		(drawing, 1419, 344, 3900, 800, 0),
		(drawing, 1420, 344, 3900, 800, 0),
		(drawing, 1421, 344, 3900, 800, 0),
		(drawing, 1422, 344, 3900, 800, 0),
		(drawing, 1423, 344, 3900, 800, 0),
		(drawing, 1424, 345, 3900, 800, 0),
		(drawing, 1425, 345, 3900, 800, 0),
		(drawing, 1426, 345, 3900, 800, 0),
		(drawing, 1427, 345, 3900, 800, 0),
		(drawing, 1428, 345, 3900, 800, 0),
		(drawing, 1429, 345, 3900, 800, 0),
		(drawing, 1430, 346, 3900, 800, 0),
		(drawing, 1431, 346, 3900, 800, 0),
		(drawing, 1432, 346, 3900, 800, 0),
		(drawing, 1433, 346, 3900, 800, 0),
		(drawing, 1434, 346, 3900, 800, 0),
		(drawing, 1435, 347, 3900, 800, 0),
		(drawing, 1436, 347, 3900, 800, 0),
		(drawing, 1437, 347, 3900, 800, 0),
		(drawing, 1438, 347, 3900, 800, 0),
		(drawing, 1439, 347, 3900, 800, 0),
		(drawing, 1440, 347, 3900, 800, 0),
		(drawing, 1441, 348, 3900, 800, 0),
		(drawing, 1442, 348, 3900, 800, 0),
		(drawing, 1443, 348, 3900, 800, 0),
		(drawing, 1444, 348, 3900, 800, 0),
		(drawing, 1445, 348, 3900, 800, 0),
		(drawing, 1446, 349, 3900, 800, 0),
		(drawing, 1447, 349, 3900, 800, 0),
		(drawing, 1448, 349, 3900, 800, 0),
		(drawing, 1449, 349, 3900, 800, 0),
		(drawing, 1450, 349, 3900, 800, 0),
		(drawing, 1451, 349, 3900, 800, 0),
		(drawing, 1452, 350, 3900, 800, 0),
		(drawing, 1453, 350, 3900, 800, 0),
		(drawing, 1454, 350, 3900, 800, 0),
		(drawing, 1455, 350, 3900, 800, 0),
		(drawing, 1456, 350, 3900, 800, 0),
		(drawing, 1457, 351, 3900, 800, 0),
		(drawing, 1458, 351, 3900, 800, 0),
		(drawing, 1459, 351, 3900, 800, 0),
		(drawing, 1460, 351, 3900, 800, 0),
		(drawing, 1461, 351, 3900, 800, 0),
		(drawing, 1462, 352, 3900, 800, 0),
		(drawing, 1463, 352, 3900, 800, 0),
		(drawing, 1464, 352, 3900, 800, 0),
		(drawing, 1465, 352, 3900, 800, 0),
		(drawing, 1466, 352, 3900, 800, 0),
		(drawing, 1467, 352, 3900, 800, 0),
		(drawing, 1468, 353, 3900, 800, 0),
		(drawing, 1469, 353, 3900, 800, 0),
		(drawing, 1470, 353, 3900, 800, 0),
		(drawing, 1471, 353, 3900, 800, 0),
		(drawing, 1472, 353, 3900, 800, 0),
		(drawing, 1473, 354, 3900, 800, 0),
		(drawing, 1474, 354, 3900, 800, 0),
		(drawing, 1475, 354, 3900, 800, 0),
		(drawing, 1476, 354, 3900, 800, 0),
		(drawing, 1477, 354, 3900, 800, 0),
		(drawing, 1478, 354, 3900, 800, 0),
		(drawing, 1479, 355, 3900, 800, 0),
		(drawing, 1480, 355, 3900, 800, 0),
		(drawing, 1481, 355, 3900, 800, 0),
		(drawing, 1482, 355, 3900, 800, 0),
		(drawing, 1483, 355, 3900, 800, 0),
		(drawing, 1484, 356, 3900, 800, 0),
		(drawing, 1485, 356, 3900, 800, 0),
		(drawing, 1486, 356, 3900, 800, 0),
		(drawing, 1487, 356, 3900, 800, 0),
		(drawing, 1488, 356, 3900, 800, 0),
		(drawing, 1489, 356, 3900, 800, 0),
		(drawing, 1490, 357, 3900, 800, 0),
		(drawing, 1491, 357, 3900, 800, 0),
		(drawing, 1492, 357, 3900, 800, 0),
		(drawing, 1493, 357, 3900, 800, 0),
		(drawing, 1494, 357, 3900, 800, 0),
		(drawing, 1495, 358, 3900, 800, 0),
		(drawing, 1496, 358, 3900, 800, 0),
		(drawing, 1497, 358, 3900, 800, 0),
		(drawing, 1498, 358, 3900, 800, 0),
		(drawing, 1499, 358, 3900, 800, 0),
		(drawing, 1500, 358, 3900, 800, 0),
		(drawing, 1501, 359, 3900, 800, 0),
		(drawing, 1502, 359, 3900, 800, 0),
		(drawing, 1503, 359, 3900, 800, 0),
		(drawing, 1504, 359, 3900, 800, 0),
		(drawing, 1505, 359, 3900, 800, 0),
		(drawing, 1506, 360, 3900, 800, 0),
		(drawing, 1507, 360, 3900, 800, 0),
		(drawing, 1508, 360, 3900, 800, 0),
		(drawing, 1509, 360, 3900, 800, 0),
		(drawing, 1510, 360, 3900, 800, 0),
		(drawing, 1511, 361, 3900, 800, 0),
		(drawing, 1512, 361, 3900, 800, 0),
		(drawing, 1513, 361, 3900, 800, 0),
		(drawing, 1514, 361, 3900, 800, 0),
		(drawing, 1515, 361, 3900, 800, 0),
		(drawing, 1516, 361, 3900, 800, 0),
		(drawing, 1517, 362, 3900, 800, 0),
		(drawing, 1518, 362, 3900, 800, 0),
		(drawing, 1519, 362, 3900, 800, 0),
		(drawing, 1520, 362, 3900, 800, 0),
		(drawing, 1521, 362, 3900, 800, 0),
		(drawing, 1522, 363, 3900, 800, 0),
		(drawing, 1523, 363, 3900, 800, 0),
		(drawing, 1524, 363, 3900, 800, 0),
		(drawing, 1525, 363, 3900, 800, 0),
		(drawing, 1526, 363, 3900, 800, 0),
		(drawing, 1527, 363, 3900, 800, 0),
		(drawing, 1528, 364, 3900, 800, 0),
		(drawing, 1529, 364, 3900, 800, 0),
		(drawing, 1530, 364, 3900, 800, 0),
		(drawing, 1531, 364, 3900, 800, 0),
		(drawing, 1532, 364, 3900, 800, 0),
		(drawing, 1533, 365, 3900, 800, 0),
		(drawing, 1534, 365, 3900, 800, 0),
		(drawing, 1535, 365, 3900, 800, 0),
		(drawing, 1536, 365, 3900, 800, 0),
		(drawing, 1537, 365, 3900, 800, 0),
		(drawing, 1538, 365, 3900, 800, 0),
		(drawing, 1539, 366, 3900, 800, 0),
		(drawing, 1540, 366, 3900, 800, 0),
		(drawing, 1541, 366, 3900, 800, 0),
		(drawing, 1542, 366, 3900, 800, 0),
		(drawing, 1543, 366, 3900, 800, 0),
		(drawing, 1544, 367, 3900, 800, 0),
		(drawing, 1545, 367, 3900, 800, 0),
		(drawing, 1546, 367, 3900, 800, 0),
		(drawing, 1547, 367, 3900, 800, 0),
		(drawing, 1548, 367, 3900, 800, 0),
		(drawing, 1549, 368, 3900, 800, 0),
		(drawing, 1550, 368, 3900, 800, 0),
		(drawing, 1551, 368, 3900, 800, 0),
		(drawing, 1552, 368, 3900, 800, 0),
		(drawing, 1553, 368, 3900, 800, 0),
		(drawing, 1554, 368, 3900, 800, 0),
		(drawing, 1555, 369, 3900, 800, 0),
		(drawing, 1556, 369, 3900, 800, 0),
		(drawing, 1557, 369, 3900, 800, 0),
		(drawing, 1558, 369, 3900, 800, 0),
		(drawing, 1559, 369, 3900, 800, 0),
		(drawing, 1560, 370, 3900, 800, 0),
		(drawing, 1561, 370, 3900, 800, 0),
		(drawing, 1562, 370, 3900, 800, 0),
		(drawing, 1563, 370, 3900, 800, 0),
		(drawing, 1564, 370, 3900, 800, 0),
		(drawing, 1565, 370, 3900, 800, 0),
		(drawing, 1566, 371, 3900, 800, 0),
		(drawing, 1567, 371, 3900, 800, 0),
		(drawing, 1568, 371, 3900, 800, 0),
		(drawing, 1569, 371, 3900, 800, 0),
		(drawing, 1570, 371, 3900, 800, 0),
		(drawing, 1571, 372, 3900, 800, 0),
		(drawing, 1572, 372, 3900, 800, 0),
		(drawing, 1573, 372, 3900, 800, 0),
		(drawing, 1574, 372, 3900, 800, 0),
		(drawing, 1575, 372, 3900, 800, 0),
		(drawing, 1576, 372, 3900, 800, 0),
		(drawing, 1577, 373, 3900, 800, 0),
		(drawing, 1578, 373, 3900, 800, 0),
		(drawing, 1579, 373, 3900, 800, 0),
		(drawing, 1580, 373, 3900, 800, 0),
		(drawing, 1581, 373, 3900, 800, 0),
		(drawing, 1582, 374, 3900, 800, 0),
		(drawing, 1583, 374, 3900, 800, 0),
		(drawing, 1584, 374, 3900, 800, 0),
		(drawing, 1585, 374, 3900, 800, 0),
		(drawing, 1586, 374, 3900, 800, 0),
		(drawing, 1587, 375, 3900, 800, 0),
		(drawing, 1588, 375, 3900, 800, 0),
		(drawing, 1589, 375, 3900, 800, 0),
		(drawing, 1590, 375, 3900, 800, 0),
		(drawing, 1591, 375, 3900, 800, 0),
		(drawing, 1592, 375, 3900, 800, 0),
		(drawing, 1593, 376, 3900, 800, 0),
		(drawing, 1594, 376, 3900, 800, 0),
		(drawing, 1595, 376, 3900, 800, 0),
		(drawing, 1596, 376, 3900, 800, 0),
		(drawing, 1597, 376, 3900, 800, 0),
		(drawing, 1598, 377, 3900, 800, 0),
		(drawing, 1599, 377, 3900, 800, 0),
		(drawing, 1600, 377, 3900, 800, 0),
		(drawing, 1601, 377, 3900, 800, 0),
		(drawing, 1602, 377, 3900, 800, 0),
		(drawing, 1603, 377, 3900, 800, 0),
		(drawing, 1604, 378, 3900, 800, 0),
		(drawing, 1605, 378, 3900, 800, 0),
		(drawing, 1606, 378, 3900, 800, 0),
		(drawing, 1607, 378, 3900, 800, 0),
		(drawing, 1608, 378, 3900, 800, 0),
		(drawing, 1609, 379, 3900, 800, 0),
		(drawing, 1610, 379, 3900, 800, 0),
		(drawing, 1611, 379, 3900, 800, 0),
		(drawing, 1612, 379, 3900, 800, 0),
		(drawing, 1613, 379, 3900, 800, 0),
		(drawing, 1614, 379, 3900, 800, 0),
		(drawing, 1615, 380, 3900, 800, 0),
		(drawing, 1616, 380, 3900, 800, 0),
		(drawing, 1617, 380, 3900, 800, 0),
		(drawing, 1618, 380, 3900, 800, 0),
		(drawing, 1619, 380, 3900, 800, 0),
		(drawing, 1620, 381, 3900, 800, 0),
		(drawing, 1621, 381, 3900, 800, 0),
		(drawing, 1622, 381, 3900, 800, 0),
		(drawing, 1623, 381, 3900, 800, 0),
		(drawing, 1624, 381, 3900, 800, 0),
		(drawing, 1625, 381, 3900, 800, 0),
		(drawing, 1626, 382, 3900, 800, 0),
		(drawing, 1627, 382, 3900, 800, 0),
		(drawing, 1628, 382, 3900, 800, 0),
		(drawing, 1629, 382, 3900, 800, 0),
		(drawing, 1630, 382, 3900, 800, 0),
		(drawing, 1631, 383, 3900, 800, 0),
		(drawing, 1632, 383, 3900, 800, 0),
		(drawing, 1633, 383, 3900, 800, 0),
		(drawing, 1634, 383, 3900, 800, 0),
		(drawing, 1635, 383, 3900, 800, 0),
		(drawing, 1636, 384, 3900, 800, 0),
		(drawing, 1637, 384, 3900, 800, 0),
		(drawing, 1638, 384, 3900, 800, 0),
		(drawing, 1639, 384, 3900, 800, 0),
		(drawing, 1640, 384, 3900, 800, 0),
		(drawing, 1641, 384, 3900, 800, 0),
		(drawing, 1642, 385, 3900, 800, 0),
		(drawing, 1643, 385, 3900, 800, 0),
		(drawing, 1644, 385, 3900, 800, 0),
		(drawing, 1645, 385, 3900, 800, 0),
		(drawing, 1646, 385, 3900, 800, 0),
		(drawing, 1647, 386, 3900, 800, 0),
		(drawing, 1648, 386, 3900, 800, 0),
		(drawing, 1649, 386, 3900, 800, 0),
		(drawing, 1650, 386, 3900, 800, 0),
		(drawing, 1651, 386, 3900, 800, 0),
		(drawing, 1652, 386, 3900, 800, 0),
		(drawing, 1653, 387, 3900, 800, 0),
		(drawing, 1654, 387, 3900, 800, 0),
		(drawing, 1655, 387, 3900, 800, 0),
		(drawing, 1656, 387, 3900, 800, 0),
		(drawing, 1657, 387, 3900, 800, 0),
		(drawing, 1658, 388, 3900, 800, 0),
		(drawing, 1659, 388, 3900, 800, 0),
		(drawing, 1660, 388, 3900, 800, 0),
		(drawing, 1661, 388, 3900, 800, 0),
		(drawing, 1662, 388, 3900, 800, 0),
		(drawing, 1663, 388, 3900, 800, 0),
		(drawing, 1664, 389, 3900, 800, 0),
		(drawing, 1665, 389, 3900, 800, 0),
		(drawing, 1666, 389, 3900, 800, 0),
		(drawing, 1667, 389, 3900, 800, 0),
		(drawing, 1668, 389, 3900, 800, 0),
		(drawing, 1669, 390, 3900, 800, 0),
		(drawing, 1670, 390, 3900, 800, 0),
		(drawing, 1671, 390, 3900, 800, 0),
		(drawing, 1672, 390, 3900, 800, 0),
		(drawing, 1673, 390, 3900, 800, 0),
		(drawing, 1674, 391, 3900, 800, 0),
		(drawing, 1675, 391, 3900, 800, 0),
		(drawing, 1676, 391, 3900, 800, 0),
		(drawing, 1677, 391, 3900, 800, 0),
		(drawing, 1678, 391, 3900, 800, 0),
		(drawing, 1679, 391, 3900, 800, 0),
		(drawing, 1680, 392, 3900, 800, 0),
		(drawing, 1681, 392, 3900, 800, 0),
		(drawing, 1682, 392, 3900, 800, 0),
		(drawing, 1683, 392, 3900, 800, 0),
		(drawing, 1684, 392, 3900, 800, 0),
		(drawing, 1685, 393, 3900, 800, 0),
		(drawing, 1686, 393, 3900, 800, 0),
		(drawing, 1687, 393, 3900, 800, 0),
		(drawing, 1688, 393, 3900, 800, 0),
		(drawing, 1689, 393, 3900, 800, 0),
		(drawing, 1690, 393, 3900, 800, 0),
		(drawing, 1691, 394, 3900, 800, 0),
		(drawing, 1692, 394, 3900, 800, 0),
		(drawing, 1693, 394, 3900, 800, 0),
		(drawing, 1694, 394, 3900, 800, 0),
		(drawing, 1695, 394, 3900, 800, 0),
		(drawing, 1696, 395, 3900, 800, 0),
		(drawing, 1697, 395, 3900, 800, 0),
		(drawing, 1698, 395, 3900, 800, 0),
		(drawing, 1699, 395, 3900, 800, 0),
		(drawing, 1700, 395, 3900, 800, 0),
		(drawing, 1701, 395, 3900, 800, 0),
		(drawing, 1702, 396, 3900, 800, 0),
		(drawing, 1703, 396, 3900, 800, 0),
		(drawing, 1704, 396, 3900, 800, 0),
		(drawing, 1705, 396, 3900, 800, 0),
		(drawing, 1706, 396, 3900, 800, 0),
		(drawing, 1707, 397, 3900, 800, 0),
		(drawing, 1708, 397, 3900, 800, 0),
		(drawing, 1709, 397, 3900, 800, 0),
		(drawing, 1710, 397, 3900, 800, 0),
		(drawing, 1711, 397, 3900, 800, 0),
		(drawing, 1712, 397, 3900, 800, 0),
		(drawing, 1713, 398, 3900, 800, 0),
		(drawing, 1714, 398, 3900, 800, 0),
		(drawing, 1715, 398, 3900, 800, 0),
		(drawing, 1716, 398, 3900, 800, 0),
		(drawing, 1717, 398, 3900, 800, 0),
		(drawing, 1718, 399, 3900, 800, 0),
		(drawing, 1719, 399, 3900, 800, 0),
		(drawing, 1720, 399, 3900, 800, 0),
		(drawing, 1721, 399, 3900, 800, 0),
		(drawing, 1722, 399, 3900, 800, 0),
		(drawing, 1723, 400, 3900, 800, 0),
		(drawing, 1724, 400, 3900, 800, 0),
		(drawing, 1725, 400, 3900, 800, 0),
		(drawing, 1726, 400, 3900, 800, 0),
		(drawing, 1727, 400, 3900, 800, 0),
		(drawing, 1728, 400, 3900, 800, 0),
		(drawing, 1729, 401, 3900, 800, 0),
		(drawing, 1730, 401, 3900, 800, 0),
		(drawing, 1731, 401, 3900, 800, 0),
		(drawing, 1732, 401, 3900, 800, 0),
		(drawing, 1733, 401, 3900, 800, 0),
		(drawing, 1734, 402, 3900, 800, 0),
		(drawing, 1735, 402, 3900, 800, 0),
		(drawing, 1736, 402, 3900, 800, 0),
		(drawing, 1737, 402, 3900, 800, 0),
		(drawing, 1738, 402, 3900, 800, 0),
		(drawing, 1739, 402, 3900, 800, 0),
		(drawing, 1740, 403, 3900, 800, 0),
		(drawing, 1741, 403, 3900, 800, 0),
		(drawing, 1742, 403, 3900, 800, 0),
		(drawing, 1743, 403, 3900, 800, 0),
		(drawing, 1744, 403, 3900, 800, 0),
		(drawing, 1745, 404, 3900, 800, 0),
		(drawing, 1746, 404, 3900, 800, 0),
		(drawing, 1747, 404, 3900, 800, 0),
		(drawing, 1748, 404, 3900, 800, 0),
		(drawing, 1749, 404, 3900, 800, 0),
		(drawing, 1750, 404, 3900, 800, 0),
		(drawing, 1751, 405, 3900, 800, 0),
		(drawing, 1752, 405, 3900, 800, 0),
		(drawing, 1753, 405, 3900, 800, 0),
		(drawing, 1754, 405, 3900, 800, 0),
		(drawing, 1755, 405, 3900, 800, 0),
		(drawing, 1756, 406, 3900, 800, 0),
		(drawing, 1757, 406, 3900, 800, 0),
		(drawing, 1758, 406, 3900, 800, 0),
		(drawing, 1759, 406, 3900, 800, 0),
		(drawing, 1760, 406, 3900, 800, 0),
		(drawing, 1761, 407, 3900, 800, 0),
		(drawing, 1762, 407, 3900, 800, 0),
		(drawing, 1763, 407, 3900, 800, 0),
		(drawing, 1764, 407, 3900, 800, 0),
		(drawing, 1765, 407, 3900, 800, 0),
		(drawing, 1766, 407, 3900, 800, 0),
		(drawing, 1767, 408, 3900, 800, 0),
		(drawing, 1768, 408, 3900, 800, 0),
		(drawing, 1769, 408, 3900, 800, 0),
		(drawing, 1770, 408, 3900, 800, 0),
		(drawing, 1771, 408, 3900, 800, 0),
		(drawing, 1772, 409, 3900, 800, 0),
		(drawing, 1773, 409, 3900, 800, 0),
		(drawing, 1774, 409, 3900, 800, 0),
		(drawing, 1775, 409, 3900, 800, 0),
		(drawing, 1776, 409, 3900, 800, 0),
		(drawing, 1777, 409, 3900, 800, 0),
		(drawing, 1778, 410, 3900, 800, 0),
		(drawing, 1779, 410, 3900, 800, 0),
		(drawing, 1780, 410, 3900, 800, 0),
		(drawing, 1781, 410, 3900, 800, 0),
		(drawing, 1782, 410, 3900, 800, 0),
		(drawing, 1783, 411, 3900, 800, 0),
		(drawing, 1784, 411, 3900, 800, 0),
		(drawing, 1785, 411, 3900, 800, 0),
		(drawing, 1786, 411, 3900, 800, 0),
		(drawing, 1787, 411, 3900, 800, 0),
		(drawing, 1788, 411, 3900, 800, 0),
		(drawing, 1789, 412, 3900, 800, 0),
		(drawing, 1790, 412, 3900, 800, 0),
		(drawing, 1791, 412, 3900, 800, 0),
		(drawing, 1792, 412, 3900, 800, 0),
		(drawing, 1793, 412, 3900, 800, 0),
		(drawing, 1794, 413, 3900, 800, 0),
		(drawing, 1795, 413, 3900, 800, 0),
		(drawing, 1796, 413, 3900, 800, 0),
		(drawing, 1797, 413, 3900, 800, 0),
		(drawing, 1798, 413, 3900, 800, 0),
		(drawing, 1799, 414, 3900, 800, 0),
		(drawing, 1800, 414, 3900, 800, 0),
		(drawing, 1801, 414, 3900, 800, 0),
		(drawing, 1802, 414, 3900, 800, 0),
		(drawing, 1803, 414, 3900, 800, 0),
		(drawing, 1804, 414, 3900, 800, 0),
		(drawing, 1805, 415, 3900, 800, 0),
		(drawing, 1806, 415, 3900, 800, 0),
		(drawing, 1807, 415, 3900, 800, 0),
		(drawing, 1808, 415, 3900, 800, 0),
		(drawing, 1809, 415, 3900, 800, 0),
		(drawing, 1810, 416, 3900, 800, 0),
		(drawing, 1811, 416, 3900, 800, 0),
		(drawing, 1812, 416, 3900, 800, 0),
		(drawing, 1813, 416, 3900, 800, 0),
		(drawing, 1814, 416, 3900, 800, 0),
		(drawing, 1815, 416, 3900, 800, 0),
		(drawing, 1816, 417, 3900, 800, 0),
		(drawing, 1817, 417, 3900, 800, 0),
		(drawing, 1818, 417, 3900, 800, 0),
		(drawing, 1819, 417, 3900, 800, 0),
		(drawing, 1820, 417, 3900, 800, 0),
		(drawing, 1821, 418, 3900, 800, 0),
		(drawing, 1822, 418, 3900, 800, 0),
		(drawing, 1823, 418, 3900, 800, 0),
		(drawing, 1824, 418, 3900, 800, 0),
		(drawing, 1825, 418, 3900, 800, 0),
		(drawing, 1826, 418, 3900, 800, 0),
		(drawing, 1827, 419, 3900, 800, 0),
		(drawing, 1828, 419, 3900, 800, 0),
		(drawing, 1829, 419, 3900, 800, 0),
		(drawing, 1830, 419, 3900, 800, 0),
		(drawing, 1831, 419, 3900, 800, 0),
		(drawing, 1832, 420, 3900, 800, 0),
		(drawing, 1833, 420, 3900, 800, 0),
		(drawing, 1834, 420, 3900, 800, 0),
		(drawing, 1835, 420, 3900, 800, 0),
		(drawing, 1836, 420, 3900, 800, 0),
		(drawing, 1837, 420, 3900, 800, 0),
		(drawing, 1838, 421, 3900, 800, 0),
		(drawing, 1839, 421, 3900, 800, 0),
		(drawing, 1840, 421, 3900, 800, 0),
		(drawing, 1841, 421, 3900, 800, 0),
		(drawing, 1842, 421, 3900, 800, 0),
		(drawing, 1843, 422, 3900, 800, 0),
		(drawing, 1844, 422, 3900, 800, 0),
		(drawing, 1845, 422, 3900, 800, 0),
		(drawing, 1846, 422, 3900, 800, 0),
		(drawing, 1847, 422, 3900, 800, 0),
		(drawing, 1848, 423, 3900, 800, 0),
		(drawing, 1849, 423, 3900, 800, 0),
		(drawing, 1850, 423, 3900, 800, 0),
		(drawing, 1851, 423, 3900, 800, 0),
		(drawing, 1852, 423, 3900, 800, 0),
		(drawing, 1853, 423, 3900, 800, 0),
		(drawing, 1854, 424, 3900, 800, 0),
		(drawing, 1855, 424, 3900, 800, 0),
		(drawing, 1856, 424, 3900, 800, 0),
		(drawing, 1857, 424, 3900, 800, 0),
		(drawing, 1858, 424, 3900, 800, 0),
		(drawing, 1859, 425, 3900, 800, 0),
		(drawing, 1860, 425, 3900, 800, 0),
		(drawing, 1861, 425, 3900, 800, 0),
		(drawing, 1862, 425, 3900, 800, 0),
		(drawing, 1863, 425, 3900, 800, 0),
		(drawing, 1864, 425, 3900, 800, 0),
		(drawing, 1865, 426, 3900, 800, 0),
		(drawing, 1866, 426, 3900, 800, 0),
		(drawing, 1867, 426, 3900, 800, 0),
		(drawing, 1868, 426, 3900, 800, 0),
		(drawing, 1869, 426, 3900, 800, 0),
		(drawing, 1870, 427, 3900, 800, 0),
		(drawing, 1871, 427, 3900, 800, 0),
		(drawing, 1872, 427, 3900, 800, 0),
		(drawing, 1873, 427, 3900, 800, 0),
		(drawing, 1874, 427, 3900, 800, 0),
		(drawing, 1875, 427, 3900, 800, 0),
		(drawing, 1876, 428, 3900, 800, 0),
		(drawing, 1877, 428, 3900, 800, 0),
		(drawing, 1878, 428, 3900, 800, 0),
		(drawing, 1879, 428, 3900, 800, 0),
		(drawing, 1880, 428, 3900, 800, 0),
		(drawing, 1881, 429, 3900, 800, 0),
		(drawing, 1882, 429, 3900, 800, 0),
		(drawing, 1883, 429, 3900, 800, 0),
		(drawing, 1884, 429, 3900, 800, 0),
		(drawing, 1885, 429, 3900, 800, 0),
		(drawing, 1886, 430, 3900, 800, 0),
		(drawing, 1887, 430, 3900, 800, 0),
		(drawing, 1888, 430, 3900, 800, 0),
		(drawing, 1889, 430, 3900, 800, 0),
		(drawing, 1890, 430, 3900, 800, 0),
		(drawing, 1891, 430, 3900, 800, 0),
		(drawing, 1892, 431, 3900, 800, 0),
		(drawing, 1893, 431, 3900, 800, 0),
		(drawing, 1894, 431, 3900, 800, 0),
		(drawing, 1895, 431, 3900, 800, 0),
		(drawing, 1896, 431, 3900, 800, 0),
		(drawing, 1897, 432, 3900, 800, 0),
		(drawing, 1898, 432, 3900, 800, 0),
		(drawing, 1899, 432, 3900, 800, 0),
		(drawing, 1900, 432, 3900, 800, 0),
		(drawing, 1901, 432, 3900, 800, 0),
		(drawing, 1902, 432, 3900, 800, 0),
		(drawing, 1903, 433, 3900, 800, 0),
		(drawing, 1904, 433, 3900, 800, 0),
		(drawing, 1905, 433, 3900, 800, 0),
		(drawing, 1906, 433, 3900, 800, 0),
		(drawing, 1907, 433, 3900, 800, 0),
		(drawing, 1908, 434, 3900, 800, 0),
		(drawing, 1909, 434, 3900, 800, 0),
		(drawing, 1910, 434, 3900, 800, 0),
		(drawing, 1911, 434, 3900, 800, 0),
		(drawing, 1912, 434, 3900, 800, 0),
		(drawing, 1913, 434, 3900, 800, 0),
		(drawing, 1914, 435, 3900, 800, 0),
		(drawing, 1915, 435, 3900, 800, 0),
		(drawing, 1916, 435, 3900, 800, 0),
		(drawing, 1917, 435, 3900, 800, 0),
		(drawing, 1918, 435, 3900, 800, 0),
		(drawing, 1919, 436, 3900, 800, 0),
		(drawing, 1920, 436, 3900, 800, 0),
		(drawing, 1921, 436, 3900, 800, 0),
		(drawing, 1922, 436, 3900, 800, 0),
		(drawing, 1923, 436, 3900, 800, 0),
		(drawing, 1924, 436, 3900, 800, 0),
		(drawing, 1925, 437, 3900, 800, 0),
		(drawing, 1926, 437, 3900, 800, 0),
		(drawing, 1927, 437, 3900, 800, 0),
		(drawing, 1928, 437, 3900, 800, 0),
		(drawing, 1929, 437, 3900, 800, 0),
		(drawing, 1930, 438, 3900, 800, 0),
		(drawing, 1931, 438, 3900, 800, 0),
		(drawing, 1932, 438, 3900, 800, 0),
		(drawing, 1933, 438, 3900, 800, 0),
		(drawing, 1934, 438, 3900, 800, 0),
		(drawing, 1935, 439, 3900, 800, 0),
		(drawing, 1936, 439, 3900, 800, 0),
		(drawing, 1937, 439, 3900, 800, 0),
		(drawing, 1938, 439, 3900, 800, 0),
		(drawing, 1939, 439, 3900, 800, 0),
		(drawing, 1940, 439, 3900, 800, 0),
		(drawing, 1941, 440, 3900, 800, 0),
		(drawing, 1942, 440, 3900, 800, 0),
		(drawing, 1943, 440, 3900, 800, 0),
		(drawing, 1944, 440, 3900, 800, 0),
		(drawing, 1945, 440, 3900, 800, 0),
		(drawing, 1946, 441, 3900, 800, 0),
		(drawing, 1947, 441, 3900, 800, 0),
		(drawing, 1948, 441, 3900, 800, 0),
		(drawing, 1949, 441, 3900, 800, 0),
		(drawing, 1950, 441, 3900, 800, 0),
		(drawing, 1951, 441, 3900, 800, 0),
		(drawing, 1952, 442, 3900, 800, 0),
		(drawing, 1953, 442, 3900, 800, 0),
		(drawing, 1954, 442, 3900, 800, 0),
		(drawing, 1955, 442, 3900, 800, 0),
		(drawing, 1956, 442, 3900, 800, 0),
		(drawing, 1957, 443, 3900, 800, 0),
		(drawing, 1958, 443, 3900, 800, 0),
		(drawing, 1959, 443, 3900, 800, 0),
		(drawing, 1960, 443, 3900, 800, 0),
		(drawing, 1961, 443, 3900, 800, 0),
		(drawing, 1962, 443, 3900, 800, 0),
		(drawing, 1963, 444, 3900, 800, 0),
		(drawing, 1964, 444, 3900, 800, 0),
		(drawing, 1965, 444, 3900, 800, 0),
		(drawing, 1966, 444, 3900, 800, 0),
		(drawing, 1967, 444, 3900, 800, 0),
		(drawing, 1968, 445, 3900, 800, 0),
		(drawing, 1969, 445, 3900, 800, 0),
		(drawing, 1970, 445, 3900, 800, 0),
		(drawing, 1971, 445, 3900, 800, 0),
		(drawing, 1972, 445, 3900, 800, 0),
		(drawing, 1973, 446, 3900, 800, 0),
		(drawing, 1974, 446, 3900, 800, 0),
		(drawing, 1975, 446, 3900, 800, 0),
		(drawing, 1976, 446, 3900, 800, 0),
		(drawing, 1977, 446, 3900, 800, 0),
		(drawing, 1978, 446, 3900, 800, 0),
		(drawing, 1979, 447, 3900, 800, 0),
		(drawing, 1980, 447, 3900, 800, 0),
		(drawing, 1981, 447, 3900, 800, 0),
		(drawing, 1982, 447, 3900, 800, 0),
		(drawing, 1983, 447, 3900, 800, 0),
		(drawing, 1984, 448, 3900, 800, 0),
		(drawing, 1985, 448, 3900, 800, 0),
		(drawing, 1986, 448, 3900, 800, 0),
		(drawing, 1987, 448, 3900, 800, 0),
		(drawing, 1988, 448, 3900, 800, 0),
		(drawing, 1989, 448, 3900, 800, 0),
		(drawing, 1990, 449, 3900, 800, 0),
		(drawing, 1991, 449, 3900, 800, 0),
		(drawing, 1992, 449, 3900, 800, 0),
		(drawing, 1993, 449, 3900, 800, 0),
		(drawing, 1994, 449, 3900, 800, 0),
		(drawing, 1995, 450, 3900, 800, 0),
		(drawing, 1996, 450, 3900, 800, 0),
		(drawing, 1997, 450, 3900, 800, 0),
		(drawing, 1998, 450, 3900, 800, 0),
		(drawing, 1999, 450, 3900, 800, 0),
		(drawing, 2000, 450, 3900, 800, 0),
		(drawing, 2001, 451, 3900, 800, 0),
		(drawing, 2002, 451, 3900, 800, 0),
		(drawing, 2003, 451, 3900, 800, 0),
		(drawing, 2004, 451, 3900, 800, 0),
		(drawing, 2005, 451, 3900, 800, 0),
		(drawing, 2006, 452, 3900, 800, 0),
		(drawing, 2007, 452, 3900, 800, 0),
		(drawing, 2008, 452, 3900, 800, 0),
		(drawing, 2009, 452, 3900, 800, 0),
		(drawing, 2010, 452, 3900, 800, 0),
		(drawing, 2011, 453, 3900, 800, 0),
		(drawing, 2012, 453, 3900, 800, 0),
		(drawing, 2013, 453, 3900, 800, 0),
		(drawing, 2014, 453, 3900, 800, 0),
		(drawing, 2015, 453, 3900, 800, 0),
		(drawing, 2016, 453, 3900, 800, 0),
		(drawing, 2017, 454, 3900, 800, 0),
		(drawing, 2018, 454, 3900, 800, 0),
		(drawing, 2019, 454, 3900, 800, 0),
		(drawing, 2020, 454, 3900, 800, 0),
		(drawing, 2021, 454, 3900, 800, 0),
		(drawing, 2022, 455, 3900, 800, 0),
		(drawing, 2023, 455, 3900, 800, 0),
		(drawing, 2024, 455, 3900, 800, 0),
		(drawing, 2025, 455, 3900, 800, 0),
		(drawing, 2026, 455, 3900, 800, 0),
		(drawing, 2027, 455, 3900, 800, 0),
		(drawing, 2028, 456, 3900, 800, 0),
		(drawing, 2029, 456, 3900, 800, 0),
		(drawing, 2030, 456, 3900, 800, 0),
		(drawing, 2031, 456, 3900, 800, 0),
		(drawing, 2032, 456, 3900, 800, 0),
		(drawing, 2033, 457, 3900, 800, 0),
		(drawing, 2034, 457, 3900, 800, 0),
		(drawing, 2035, 457, 3900, 800, 0),
		(drawing, 2036, 457, 3900, 800, 0),
		(drawing, 2037, 457, 3900, 800, 0),
		(drawing, 2038, 457, 3900, 800, 0),
		(drawing, 2039, 458, 3900, 800, 0),
		(drawing, 2040, 458, 3900, 800, 0),
		(drawing, 2041, 458, 3900, 800, 0),
		(drawing, 2042, 458, 3900, 800, 0),
		(drawing, 2043, 458, 3900, 800, 0),
		(drawing, 2044, 459, 3900, 800, 0),
		(drawing, 2045, 459, 3900, 800, 0),
		(drawing, 2046, 459, 3900, 800, 0),
		(drawing, 2047, 459, 3900, 800, 0),
		(drawing, 2048, 459, 3900, 800, 0),
		(drawing, 2049, 459, 3900, 800, 0),
		(drawing, 2050, 460, 3900, 800, 0),
		(drawing, 2051, 460, 3900, 800, 0),
		(drawing, 2052, 460, 3900, 800, 0),
		(drawing, 2053, 460, 3900, 800, 0),
		(drawing, 2054, 460, 3900, 800, 0),
		(drawing, 2055, 461, 3900, 800, 0),
		(drawing, 2056, 461, 3900, 800, 0),
		(drawing, 2057, 461, 3900, 800, 0),
		(drawing, 2058, 461, 3900, 800, 0),
		(drawing, 2059, 461, 3900, 800, 0),
		(drawing, 2060, 462, 3900, 800, 0),
		(drawing, 2061, 462, 3900, 800, 0),
		(drawing, 2062, 462, 3900, 800, 0),
		(drawing, 2063, 462, 3900, 800, 0),
		(drawing, 2064, 462, 3900, 800, 0),
		(drawing, 2065, 462, 3900, 800, 0),
		(drawing, 2066, 463, 3900, 800, 0),
		(drawing, 2067, 463, 3900, 800, 0),
		(drawing, 2068, 463, 3900, 800, 0),
		(drawing, 2069, 463, 3900, 800, 0),
		(drawing, 2070, 463, 3900, 800, 0),
		(drawing, 2071, 464, 3900, 800, 0),
		(drawing, 2072, 464, 3900, 800, 0),
		(drawing, 2073, 464, 3900, 800, 0),
		(drawing, 2074, 464, 3900, 800, 0),
		(drawing, 2075, 464, 3900, 800, 0),
		(drawing, 2076, 464, 3900, 800, 0),
		(drawing, 2077, 465, 3900, 800, 0),
		(drawing, 2078, 465, 3900, 800, 0),
		(drawing, 2079, 465, 3900, 800, 0),
		(drawing, 2080, 465, 3900, 800, 0),
		(drawing, 2081, 465, 3900, 800, 0),
		(drawing, 2082, 466, 3900, 800, 0),
		(drawing, 2083, 466, 3900, 800, 0),
		(drawing, 2084, 466, 3900, 800, 0),
		(drawing, 2085, 466, 3900, 800, 0),
		(drawing, 2086, 466, 3900, 800, 0),
		(drawing, 2087, 466, 3900, 800, 0),
		(drawing, 2088, 467, 3900, 800, 0),
		(drawing, 2089, 467, 3900, 800, 0),
		(drawing, 2090, 467, 3900, 800, 0),
		(drawing, 2091, 467, 3900, 800, 0),
		(drawing, 2092, 467, 3900, 800, 0),
		(drawing, 2093, 468, 3900, 800, 0),
		(drawing, 2094, 468, 3900, 800, 0),
		(drawing, 2095, 468, 3900, 800, 0),
		(drawing, 2096, 468, 3900, 800, 0),
		(drawing, 2097, 468, 3900, 800, 0),
		(drawing, 2098, 469, 3900, 800, 0),
		(drawing, 2099, 469, 3900, 800, 0),
		(drawing, 2100, 469, 3900, 800, 0),
		(drawing, 2101, 469, 3900, 800, 0),
		(drawing, 2102, 469, 3900, 800, 0),
		(drawing, 2103, 469, 3900, 800, 0),
		(drawing, 2104, 470, 3900, 800, 0),
		(drawing, 2105, 470, 3900, 800, 0),
		(drawing, 2106, 470, 3900, 800, 0),
		(drawing, 2107, 470, 3900, 800, 0),
		(drawing, 2108, 470, 3900, 800, 0),
		(drawing, 2109, 471, 3900, 800, 0),
		(drawing, 2110, 471, 3900, 800, 0),
		(drawing, 2111, 471, 3900, 800, 0),
		(drawing, 2112, 471, 3900, 800, 0),
		(drawing, 2113, 471, 3900, 800, 0),
		(drawing, 2114, 471, 3900, 800, 0),
		(drawing, 2115, 472, 3900, 800, 0),
		(drawing, 2116, 472, 3900, 800, 0),
		(drawing, 2117, 472, 3900, 800, 0),
		(drawing, 2118, 472, 3900, 800, 0),
		(drawing, 2119, 472, 3900, 800, 0),
		(drawing, 2120, 473, 3900, 800, 0),
		(drawing, 2121, 473, 3900, 800, 0),
		(drawing, 2122, 473, 3900, 800, 0),
		(drawing, 2123, 473, 3900, 800, 0),
		(drawing, 2124, 473, 3900, 800, 0),
		(drawing, 2125, 473, 3900, 800, 0),
		(drawing, 2126, 474, 3900, 800, 0),
		(drawing, 2127, 474, 3900, 800, 0),
		(drawing, 2128, 474, 3900, 800, 0),
		(drawing, 2129, 474, 3900, 800, 0),
		(drawing, 2130, 474, 3900, 800, 0),
		(drawing, 2131, 475, 3900, 800, 0),
		(drawing, 2132, 475, 3900, 800, 0),
		(drawing, 2133, 475, 3900, 800, 0),
		(drawing, 2134, 475, 3900, 800, 0),
		(drawing, 2135, 475, 3900, 800, 0),
		(drawing, 2136, 475, 3900, 800, 0),
		(drawing, 2137, 476, 3900, 800, 0),
		(drawing, 2138, 476, 3900, 800, 0),
		(drawing, 2139, 476, 3900, 800, 0),
		(drawing, 2140, 476, 3900, 800, 0),
		(drawing, 2141, 476, 3900, 800, 0),
		(drawing, 2142, 477, 3900, 800, 0),
		(drawing, 2143, 477, 3900, 800, 0),
		(drawing, 2144, 477, 3900, 800, 0),
		(drawing, 2145, 477, 3900, 800, 0),
		(drawing, 2146, 477, 3900, 800, 0),
		(drawing, 2147, 478, 3900, 800, 0),
		(drawing, 2148, 478, 3900, 800, 0),
		(drawing, 2149, 478, 3900, 800, 0),
		(drawing, 2150, 478, 3900, 800, 0),
		(drawing, 2151, 478, 3900, 800, 0),
		(drawing, 2152, 478, 3900, 800, 0),
		(drawing, 2153, 479, 3900, 800, 0),
		(drawing, 2154, 479, 3900, 800, 0),
		(drawing, 2155, 479, 3900, 800, 0),
		(drawing, 2156, 479, 3900, 800, 0),
		(drawing, 2157, 479, 3900, 800, 0),
		(drawing, 2158, 480, 3900, 800, 0),
		(drawing, 2159, 480, 3900, 800, 0),
		(drawing, 2160, 480, 3900, 800, 0),
		(drawing, 2161, 480, 3900, 800, 0),
		(drawing, 2162, 480, 3900, 800, 0),
		(drawing, 2163, 480, 3900, 800, 0),
		(drawing, 2164, 481, 3900, 800, 0),
		(drawing, 2165, 481, 3900, 800, 0),
		(drawing, 2166, 481, 3900, 800, 0),
		(drawing, 2167, 481, 3900, 800, 0),
		(drawing, 2168, 481, 3900, 800, 0),
		(drawing, 2169, 482, 3900, 800, 0),
		(drawing, 2170, 482, 3900, 800, 0),
		(drawing, 2171, 482, 3900, 800, 0),
		(drawing, 2172, 482, 3900, 800, 0),
		(drawing, 2173, 482, 3900, 800, 0),
		(drawing, 2174, 482, 3900, 800, 0),
		(drawing, 2175, 483, 3900, 800, 0),
		(drawing, 2176, 483, 3900, 800, 0),
		(drawing, 2177, 483, 3900, 800, 0),
		(drawing, 2178, 483, 3900, 800, 0),
		(drawing, 2179, 483, 3900, 800, 0),
		(drawing, 2180, 484, 3900, 800, 0),
		(drawing, 2181, 484, 3900, 800, 0),
		(drawing, 2182, 484, 3900, 800, 0),
		(drawing, 2183, 484, 3900, 800, 0),
		(drawing, 2184, 484, 3900, 800, 0),
		(drawing, 2185, 485, 3900, 800, 0),
		(drawing, 2186, 485, 3900, 800, 0),
		(drawing, 2187, 485, 3900, 800, 0),
		(drawing, 2188, 485, 3900, 800, 0),
		(drawing, 2189, 485, 3900, 800, 0),
		(drawing, 2190, 485, 3900, 800, 0),
		(drawing, 2191, 486, 3900, 800, 0),
		(drawing, 2192, 486, 3900, 800, 0),
		(drawing, 2193, 486, 3900, 800, 0),
		(drawing, 2194, 486, 3900, 800, 0),
		(drawing, 2195, 486, 3900, 800, 0),
		(drawing, 2196, 487, 3900, 800, 0),
		(drawing, 2197, 487, 3900, 800, 0),
		(drawing, 2198, 487, 3900, 800, 0),
		(drawing, 2199, 487, 3900, 800, 0),
		(drawing, 2200, 487, 3900, 800, 0),
		(drawing, 2201, 487, 3900, 800, 0),
		(drawing, 2202, 488, 3900, 800, 0),
		(drawing, 2203, 488, 3900, 800, 0),
		(drawing, 2204, 488, 3900, 800, 0),
		(drawing, 2205, 488, 3900, 800, 0),
		(drawing, 2206, 488, 3900, 800, 0),
		(drawing, 2207, 489, 3900, 800, 0),
		(drawing, 2208, 489, 3900, 800, 0),
		(drawing, 2209, 489, 3900, 800, 0),
		(drawing, 2210, 489, 3900, 800, 0),
		(drawing, 2211, 489, 3900, 800, 0),
		(drawing, 2212, 489, 3900, 800, 0),
		(drawing, 2213, 490, 3900, 800, 0),
		(drawing, 2214, 490, 3900, 800, 0),
		(drawing, 2215, 490, 3900, 800, 0),
		(drawing, 2216, 490, 3900, 800, 0),
		(drawing, 2217, 490, 3900, 800, 0),
		(drawing, 2218, 491, 3900, 800, 0),
		(drawing, 2219, 491, 3900, 800, 0),
		(drawing, 2220, 491, 3900, 800, 0),
		(drawing, 2221, 491, 3900, 800, 0),
		(drawing, 2222, 491, 3900, 800, 0),
		(drawing, 2223, 492, 3900, 800, 0),
		(drawing, 2224, 492, 3900, 800, 0),
		(drawing, 2225, 492, 3900, 800, 0),
		(drawing, 2226, 492, 3900, 800, 0),
		(drawing, 2227, 492, 3900, 800, 0),
		(drawing, 2228, 492, 3900, 800, 0),
		(drawing, 2229, 493, 3900, 800, 0),
		(drawing, 2230, 493, 3900, 800, 0),
		(drawing, 2231, 493, 3900, 800, 0),
		(drawing, 2232, 493, 3900, 800, 0),
		(drawing, 2233, 493, 3900, 800, 0),
		(drawing, 2234, 494, 3900, 800, 0),
		(drawing, 2235, 494, 3900, 800, 0),
		(drawing, 2236, 494, 3900, 800, 0),
		(drawing, 2237, 494, 3900, 800, 0),
		(drawing, 2238, 494, 3900, 800, 0),
		(drawing, 2239, 494, 3900, 800, 0),
		(drawing, 2240, 495, 3900, 800, 0),
		(drawing, 2241, 495, 3900, 800, 0),
		(drawing, 2242, 495, 3900, 800, 0),
		(drawing, 2243, 495, 3900, 800, 0),
		(drawing, 2244, 495, 3900, 800, 0),
		(drawing, 2245, 496, 3900, 800, 0),
		(drawing, 2246, 496, 3900, 800, 0),
		(drawing, 2247, 496, 3900, 800, 0),
		(drawing, 2248, 496, 3900, 800, 0),
		(drawing, 2249, 496, 3900, 800, 0),
		(drawing, 2250, 496, 3900, 800, 0),
		(drawing, 2251, 497, 3900, 800, 0),
		(drawing, 2252, 497, 3900, 800, 0),
		(drawing, 2253, 497, 3900, 800, 0),
		(drawing, 2254, 497, 3900, 800, 0),
		(drawing, 2255, 497, 3900, 800, 0),
		(drawing, 2256, 498, 3900, 800, 0),
		(drawing, 2257, 498, 3900, 800, 0),
		(drawing, 2258, 498, 3900, 800, 0),
		(drawing, 2259, 498, 3900, 800, 0),
		(drawing, 2260, 498, 3900, 800, 0),
		(drawing, 2261, 498, 3900, 800, 0),
		(drawing, 2262, 499, 3900, 800, 0),
		(drawing, 2263, 499, 3900, 800, 0),
		(drawing, 2264, 499, 3900, 800, 0),
		(drawing, 2265, 499, 3900, 800, 0),
		(drawing, 2266, 499, 3900, 800, 0),
		(drawing, 2267, 500, 3900, 800, 0),
		(drawing, 2268, 500, 3900, 800, 0),
		(drawing, 2269, 500, 3900, 800, 0),
		(drawing, 2270, 500, 3900, 800, 0),
		(drawing, 2271, 500, 3900, 800, 0),
		(drawing, 2272, 501, 3900, 800, 0),
		(drawing, 2273, 501, 3900, 800, 0),
		(drawing, 2274, 501, 3900, 800, 0),
		(drawing, 2275, 501, 3900, 800, 0),
		(drawing, 2276, 501, 3900, 800, 0),
		(drawing, 2277, 501, 3900, 800, 0),
		(drawing, 2278, 502, 3900, 800, 0),
		(drawing, 2279, 502, 3900, 800, 0),
		(drawing, 2280, 502, 3900, 800, 0),
		(drawing, 2281, 502, 3900, 800, 0),
		(drawing, 2282, 502, 3900, 800, 0),
		(drawing, 2283, 503, 3900, 800, 0),
		(drawing, 2284, 503, 3900, 800, 0),
		(drawing, 2285, 503, 3900, 800, 0),
		(drawing, 2286, 503, 3900, 800, 0),
		(drawing, 2287, 503, 3900, 800, 0),
		(drawing, 2288, 503, 3900, 800, 0),
		(drawing, 2289, 504, 3900, 800, 0),
		(drawing, 2290, 504, 3900, 800, 0),
		(drawing, 2291, 504, 3900, 800, 0),
		(drawing, 2292, 504, 3900, 800, 0),
		(drawing, 2293, 504, 3900, 800, 0),
		(drawing, 2294, 505, 3900, 800, 0),
		(drawing, 2295, 505, 3900, 800, 0),
		(drawing, 2296, 505, 3900, 800, 0),
		(drawing, 2297, 505, 3900, 800, 0),
		(drawing, 2298, 505, 3900, 800, 0),
		(drawing, 2299, 505, 3900, 800, 0),
		(drawing, 2300, 506, 3900, 800, 0),
		(drawing, 2301, 506, 3900, 800, 0),
		(drawing, 2302, 506, 3900, 800, 0),
		(drawing, 2303, 506, 3900, 800, 0),
		(drawing, 2304, 506, 3900, 800, 0),
		(drawing, 2305, 507, 3900, 800, 0),
		(drawing, 2306, 507, 3900, 800, 0),
		(drawing, 2307, 507, 3900, 800, 0),
		(drawing, 2308, 507, 3900, 800, 0),
		(drawing, 2309, 507, 3900, 800, 0),
		(drawing, 2310, 508, 3900, 800, 0),
		(drawing, 2311, 508, 3900, 800, 0),
		(drawing, 2312, 508, 3900, 800, 0),
		(drawing, 2313, 508, 3900, 800, 0),
		(drawing, 2314, 508, 3900, 800, 0),
		(drawing, 2315, 508, 3900, 800, 0),
		(drawing, 2316, 509, 3900, 800, 0),
		(drawing, 2317, 509, 3900, 800, 0),
		(drawing, 2318, 509, 3900, 800, 0),
		(drawing, 2319, 509, 3900, 800, 0),
		(drawing, 2320, 509, 3900, 800, 0),
		(drawing, 2321, 510, 3900, 800, 0),
		(drawing, 2322, 510, 3900, 800, 0),
		(drawing, 2323, 510, 3900, 800, 0),
		(drawing, 2324, 510, 3900, 800, 0),
		(drawing, 2325, 510, 3900, 800, 0),
		(drawing, 2326, 510, 3900, 800, 0),
		(drawing, 2327, 511, 3900, 800, 0),
		(drawing, 2328, 511, 3900, 800, 0),
		(drawing, 2329, 511, 3900, 800, 0),
		(drawing, 2330, 511, 3900, 800, 0),
		(drawing, 2331, 511, 3900, 800, 0),
		(drawing, 2332, 512, 3900, 800, 0),
		(drawing, 2333, 512, 3900, 800, 0),
		(drawing, 2334, 512, 3900, 800, 0),
		(drawing, 2335, 512, 3900, 800, 0),
		(drawing, 2336, 512, 3900, 800, 0),
		(drawing, 2337, 512, 3900, 800, 0),
		(drawing, 2338, 513, 3900, 800, 0),
		(drawing, 2339, 513, 3900, 800, 0),
		(drawing, 2340, 513, 3900, 800, 0),
		(drawing, 2341, 513, 3900, 800, 0),
		(drawing, 2342, 513, 3900, 800, 0),
		(drawing, 2343, 514, 3900, 800, 0),
		(drawing, 2344, 514, 3900, 800, 0),
		(drawing, 2345, 514, 3900, 800, 0),
		(drawing, 2346, 514, 3900, 800, 0),
		(drawing, 2347, 514, 3900, 800, 0),
		(drawing, 2348, 514, 3900, 800, 0),
		(drawing, 2349, 515, 3900, 800, 0),
		(drawing, 2350, 515, 3900, 800, 0),
		(drawing, 2351, 515, 3900, 800, 0),
		(drawing, 2352, 515, 3900, 800, 0),
		(drawing, 2353, 515, 3900, 800, 0),
		(drawing, 2354, 516, 3900, 800, 0),
		(drawing, 2355, 516, 3900, 800, 0),
		(drawing, 2356, 516, 3900, 800, 0),
		(drawing, 2357, 516, 3900, 800, 0),
		(drawing, 2358, 516, 3900, 800, 0),
		(drawing, 2359, 517, 3900, 800, 0),
		(drawing, 2360, 517, 3900, 800, 0),
		(drawing, 2361, 517, 3900, 800, 0),
		(drawing, 2362, 517, 3900, 800, 0),
		(drawing, 2363, 517, 3900, 800, 0),
		(drawing, 2364, 517, 3900, 800, 0),
		(drawing, 2365, 518, 3900, 800, 0),
		(drawing, 2366, 518, 3900, 800, 0),
		(drawing, 2367, 518, 3900, 800, 0),
		(drawing, 2368, 518, 3900, 800, 0),
		(drawing, 2369, 518, 3900, 800, 0),
		(drawing, 2370, 519, 3900, 800, 0),
		(drawing, 2371, 519, 3900, 800, 0),
		(drawing, 2372, 519, 3900, 800, 0),
		(drawing, 2373, 519, 3900, 800, 0),
		(drawing, 2374, 519, 3900, 800, 0),
		(drawing, 2375, 519, 3900, 800, 0),
		(drawing, 2376, 520, 3900, 800, 0),
		(drawing, 2377, 520, 3900, 800, 0),
		(drawing, 2378, 520, 3900, 800, 0),
		(drawing, 2379, 520, 3900, 800, 0),
		(drawing, 2380, 520, 3900, 800, 0),
		(drawing, 2381, 521, 3900, 800, 0),
		(drawing, 2382, 521, 3900, 800, 0),
		(drawing, 2383, 521, 3900, 800, 0),
		(drawing, 2384, 521, 3900, 800, 0),
		(drawing, 2385, 521, 3900, 800, 0),
		(drawing, 2386, 521, 3900, 800, 0),
		(drawing, 2387, 522, 3900, 800, 0),
		(drawing, 2388, 522, 3900, 800, 0),
		(drawing, 2389, 522, 3900, 800, 0),
		(drawing, 2390, 522, 3900, 800, 0),
		(drawing, 2391, 522, 3900, 800, 0),
		(drawing, 2392, 523, 3900, 800, 0),
		(drawing, 2393, 523, 3900, 800, 0),
		(drawing, 2394, 523, 3900, 800, 0),
		(drawing, 2395, 523, 3900, 800, 0),
		(drawing, 2396, 523, 3900, 800, 0),
		(drawing, 2397, 524, 3900, 800, 0),
		(drawing, 2398, 524, 3900, 800, 0),
		(drawing, 2399, 524, 3900, 800, 0),
		(drawing, 2400, 524, 3900, 800, 0),
		(drawing, 2401, 524, 3900, 800, 0),
		(drawing, 2402, 524, 3900, 800, 0),
		(drawing, 2403, 525, 3900, 800, 0),
		(drawing, 2404, 525, 3900, 800, 0),
		(drawing, 2405, 525, 3900, 800, 0),
		(drawing, 2406, 525, 3900, 800, 0),
		(drawing, 2407, 525, 3900, 800, 0),
		(drawing, 2408, 526, 3900, 800, 0),
		(drawing, 2409, 526, 3900, 800, 0),
		(drawing, 2410, 526, 3900, 800, 0),
		(drawing, 2411, 526, 3900, 800, 0),
		(drawing, 2412, 526, 3900, 800, 0),
		(drawing, 2413, 526, 3900, 800, 0),
		(drawing, 2414, 527, 3900, 800, 0),
		(drawing, 2415, 527, 3900, 800, 0),
		(drawing, 2416, 527, 3900, 800, 0),
		(drawing, 2417, 527, 3900, 800, 0),
		(drawing, 2418, 527, 3900, 800, 0),
		(drawing, 2419, 528, 3900, 800, 0),
		(drawing, 2420, 528, 3900, 800, 0),
		(drawing, 2421, 528, 3900, 800, 0),
		(drawing, 2422, 528, 3900, 800, 0),
		(drawing, 2423, 528, 3900, 800, 0),
		(drawing, 2424, 528, 3900, 800, 0),
		(drawing, 2425, 529, 3900, 800, 0),
		(drawing, 2426, 529, 3900, 800, 0),
		(drawing, 2427, 529, 3900, 800, 0),
		(drawing, 2428, 529, 3900, 800, 0),
		(drawing, 2429, 529, 3900, 800, 0),
		(drawing, 2430, 530, 3900, 800, 0),
		(drawing, 2431, 530, 3900, 800, 0),
		(drawing, 2432, 530, 3900, 800, 0),
		(drawing, 2433, 530, 3900, 800, 0),
		(drawing, 2434, 530, 3900, 800, 0),
		(drawing, 2435, 531, 3900, 800, 0),
		(drawing, 2436, 531, 3900, 800, 0),
		(drawing, 2437, 531, 3900, 800, 0),
		(drawing, 2438, 531, 3900, 800, 0),
		(drawing, 2439, 531, 3900, 800, 0),
		(drawing, 2440, 531, 3900, 800, 0),
		(drawing, 2441, 532, 3900, 800, 0),
		(drawing, 2442, 532, 3900, 800, 0),
		(drawing, 2443, 532, 3900, 800, 0),
		(drawing, 2444, 532, 3900, 800, 0),
		(drawing, 2445, 532, 3900, 800, 0),
		(drawing, 2446, 533, 3900, 800, 0),
		(drawing, 2447, 533, 3900, 800, 0),
		(drawing, 2448, 533, 3900, 800, 0),
		(drawing, 2449, 533, 3900, 800, 0),
		(drawing, 2450, 533, 3900, 800, 0),
		(drawing, 2451, 533, 3900, 800, 0),
		(drawing, 2452, 534, 3900, 800, 0),
		(drawing, 2453, 534, 3900, 800, 0),
		(drawing, 2454, 534, 3900, 800, 0),
		(drawing, 2455, 534, 3900, 800, 0),
		(drawing, 2456, 534, 3900, 800, 0),
		(drawing, 2457, 535, 3900, 800, 0),
		(drawing, 2458, 535, 3900, 800, 0),
		(drawing, 2459, 535, 3900, 800, 0),
		(drawing, 2460, 535, 3900, 800, 0),
		(drawing, 2461, 535, 3900, 800, 0),
		(drawing, 2462, 535, 3900, 800, 0),
		(drawing, 2463, 536, 3900, 800, 0),
		(drawing, 2464, 536, 3900, 800, 0),
		(drawing, 2465, 536, 3900, 800, 0),
		(drawing, 2466, 536, 3900, 800, 0),
		(drawing, 2467, 536, 3900, 800, 0),
		(drawing, 2468, 537, 3900, 800, 0),
		(drawing, 2469, 537, 3900, 800, 0),
		(drawing, 2470, 537, 3900, 800, 0),
		(drawing, 2471, 537, 3900, 800, 0),
		(drawing, 2472, 537, 3900, 800, 0),
		(drawing, 2473, 537, 3900, 800, 0),
		(drawing, 2474, 538, 3900, 800, 0),
		(drawing, 2475, 538, 3900, 800, 0),
		(drawing, 2476, 538, 3900, 800, 0),
		(drawing, 2477, 538, 3900, 800, 0),
		(drawing, 2478, 538, 3900, 800, 0),
		(drawing, 2479, 539, 3900, 800, 0),
		(drawing, 2480, 539, 3900, 800, 0),
		(drawing, 2481, 539, 3900, 800, 0),
		(drawing, 2482, 539, 3900, 800, 0),
		(drawing, 2483, 539, 3900, 800, 0),
		(drawing, 2484, 540, 3900, 800, 0),
		(drawing, 2485, 540, 3900, 800, 0),
		(drawing, 2486, 540, 3900, 800, 0),
		(drawing, 2487, 540, 3900, 800, 0),
		(drawing, 2488, 540, 3900, 800, 0),
		(drawing, 2489, 540, 3900, 800, 0),
		(drawing, 2490, 541, 3900, 800, 0),
		(drawing, 2491, 541, 3900, 800, 0),
		(drawing, 2492, 541, 3900, 800, 0),
		(drawing, 2493, 541, 3900, 800, 0),
		(drawing, 2494, 541, 3900, 800, 0),
		(drawing, 2495, 542, 3900, 800, 0),
		(drawing, 2496, 542, 3900, 800, 0),
		(drawing, 2497, 542, 3900, 800, 0),
		(drawing, 2498, 542, 3900, 800, 0),
		(drawing, 2499, 542, 3900, 800, 0),
		(drawing, 2500, 542, 3900, 800, 0),
		(drawing, 2501, 543, 3900, 800, 0),
		(drawing, 2502, 543, 3900, 800, 0),
		(drawing, 2503, 543, 3900, 800, 0),
		(drawing, 2504, 543, 3900, 800, 0),
		(drawing, 2505, 543, 3900, 800, 0),
		(drawing, 2506, 544, 3900, 800, 0),
		(drawing, 2507, 544, 3900, 800, 0),
		(drawing, 2508, 544, 3900, 800, 0),
		(drawing, 2509, 544, 3900, 800, 0),
		(drawing, 2510, 544, 3900, 800, 0),
		(drawing, 2511, 544, 3900, 800, 0),
		(drawing, 2512, 545, 3900, 800, 0),
		(drawing, 2513, 545, 3900, 800, 0),
		(drawing, 2514, 545, 3900, 800, 0),
		(drawing, 2515, 545, 3900, 800, 0),
		(drawing, 2516, 545, 3900, 800, 0),
		(drawing, 2517, 546, 3900, 800, 0),
		(drawing, 2518, 546, 3900, 800, 0),
		(drawing, 2519, 546, 3900, 800, 0),
		(drawing, 2520, 546, 3900, 800, 0),
		(drawing, 2521, 546, 3900, 800, 0),
		(drawing, 2522, 547, 3900, 800, 0),
		(drawing, 2523, 547, 3900, 800, 0),
		(drawing, 2524, 547, 3900, 800, 0),
		(drawing, 2525, 547, 3900, 800, 0),
		(drawing, 2526, 547, 3900, 800, 0),
		(drawing, 2527, 547, 3900, 800, 0),
		(drawing, 2528, 548, 3900, 800, 0),
		(drawing, 2529, 548, 3900, 800, 0),
		(drawing, 2530, 548, 3900, 800, 0),
		(drawing, 2531, 548, 3900, 800, 0),
		(drawing, 2532, 548, 3900, 800, 0),
		(drawing, 2533, 549, 3900, 800, 0),
		(drawing, 2534, 549, 3900, 800, 0),
		(drawing, 2535, 549, 3900, 800, 0),
		(drawing, 2536, 549, 3900, 800, 0),
		(drawing, 2537, 549, 3900, 800, 0),
		(drawing, 2538, 549, 3900, 800, 0),
		(drawing, 2539, 550, 3900, 800, 0),
		(drawing, 2540, 550, 3900, 800, 0),
		(drawing, 2541, 550, 3900, 800, 0),
		(drawing, 2542, 550, 3900, 800, 0),
		(drawing, 2543, 550, 3900, 800, 0),
		(drawing, 2544, 551, 3900, 800, 0),
		(drawing, 2545, 551, 3900, 800, 0),
		(drawing, 2546, 551, 3900, 800, 0),
		(drawing, 2547, 551, 3900, 800, 0),
		(drawing, 2548, 551, 3900, 800, 0),
		(drawing, 2549, 551, 3900, 800, 0),
		(drawing, 2550, 552, 3900, 800, 0),
		(drawing, 2551, 552, 3900, 800, 0),
		(drawing, 2552, 552, 3900, 800, 0),
		(drawing, 2553, 552, 3900, 800, 0),
		(drawing, 2554, 552, 3900, 800, 0),
		(drawing, 2555, 553, 3900, 800, 0),
		(drawing, 2556, 553, 3900, 800, 0),
		(drawing, 2557, 553, 3900, 800, 0),
		(drawing, 2558, 553, 3900, 800, 0),
		(drawing, 2559, 553, 3900, 800, 0),
		(drawing, 2560, 553, 3900, 800, 0),
		(drawing, 2561, 554, 3900, 800, 0),
		(drawing, 2562, 554, 3900, 800, 0),
		(drawing, 2563, 554, 3900, 800, 0),
		(drawing, 2564, 554, 3900, 800, 0),
		(drawing, 2565, 554, 3900, 800, 0),
		(drawing, 2566, 555, 3900, 800, 0),
		(drawing, 2567, 555, 3900, 800, 0),
		(drawing, 2568, 555, 3900, 800, 0),
		(drawing, 2569, 555, 3900, 800, 0),
		(drawing, 2570, 555, 3900, 800, 0),
		(drawing, 2571, 556, 3900, 800, 0),
		(drawing, 2572, 556, 3900, 800, 0),
		(drawing, 2573, 556, 3900, 800, 0),
		(drawing, 2574, 556, 3900, 800, 0),
		(drawing, 2575, 556, 3900, 800, 0),
		(drawing, 2576, 556, 3900, 800, 0),
		(drawing, 2577, 557, 3900, 800, 0),
		(drawing, 2578, 557, 3900, 800, 0),
		(drawing, 2579, 557, 3900, 800, 0),
		(drawing, 2580, 557, 3900, 800, 0),
		(drawing, 2581, 557, 3900, 800, 0),
		(drawing, 2582, 558, 3900, 800, 0),
		(drawing, 2583, 558, 3900, 800, 0),
		(drawing, 2584, 558, 3900, 800, 0),
		(drawing, 2585, 558, 3900, 800, 0),
		(drawing, 2586, 558, 3900, 800, 0),
		(drawing, 2587, 558, 3900, 800, 0),
		(drawing, 2588, 559, 3900, 800, 0),
		(drawing, 2589, 559, 3900, 800, 0),
		(drawing, 2590, 559, 3900, 800, 0),
		(drawing, 2591, 559, 3900, 800, 0),
		(drawing, 2592, 559, 3900, 800, 0),
		(drawing, 2593, 560, 3900, 800, 0),
		(drawing, 2594, 560, 3900, 800, 0),
		(drawing, 2595, 560, 3900, 800, 0),
		(drawing, 2596, 560, 3900, 800, 0),
		(drawing, 2597, 560, 3900, 800, 0),
		(drawing, 2598, 560, 3900, 800, 0),
		(drawing, 2599, 561, 3900, 800, 0),
		(drawing, 2600, 561, 3900, 800, 0),
		(drawing, 2601, 561, 3900, 800, 0),
		(drawing, 2602, 561, 3900, 800, 0),
		(drawing, 2603, 561, 3900, 800, 0),
		(drawing, 2604, 562, 3900, 800, 0),
		(drawing, 2605, 562, 3900, 800, 0),
		(drawing, 2606, 562, 3900, 800, 0),
		(drawing, 2607, 562, 3900, 800, 0),
		(drawing, 2608, 562, 3900, 800, 0),
		(drawing, 2609, 563, 3900, 800, 0),
		(drawing, 2610, 563, 3900, 800, 0),
		(drawing, 2611, 563, 3900, 800, 0),
		(drawing, 2612, 563, 3900, 800, 0),
		(drawing, 2613, 563, 3900, 800, 0),
		(drawing, 2614, 563, 3900, 800, 0),
		(drawing, 2615, 564, 3900, 800, 0),
		(drawing, 2616, 564, 3900, 800, 0),
		(drawing, 2617, 564, 3900, 800, 0),
		(drawing, 2618, 564, 3900, 800, 0),
		(drawing, 2619, 564, 3900, 800, 0),
		(drawing, 2620, 565, 3900, 800, 0),
		(drawing, 2621, 565, 3900, 800, 0),
		(drawing, 2622, 565, 3900, 800, 0),
		(drawing, 2623, 565, 3900, 800, 0),
		(drawing, 2624, 565, 3900, 800, 0),
		(drawing, 2625, 565, 3900, 800, 0),
		(drawing, 2626, 566, 3900, 800, 0),
		(drawing, 2627, 566, 3900, 800, 0),
		(drawing, 2628, 566, 3900, 800, 0),
		(drawing, 2629, 566, 3900, 800, 0),
		(drawing, 2630, 566, 3900, 800, 0),
		(drawing, 2631, 567, 3900, 800, 0),
		(drawing, 2632, 567, 3900, 800, 0),
		(drawing, 2633, 567, 3900, 800, 0),
		(drawing, 2634, 567, 3900, 800, 0),
		(drawing, 2635, 567, 3900, 800, 0),
		(drawing, 2636, 567, 3900, 800, 0),
		(drawing, 2637, 568, 3900, 800, 0),
		(drawing, 2638, 568, 3900, 800, 0),
		(drawing, 2639, 568, 3900, 800, 0),
		(drawing, 2640, 568, 3900, 800, 0),
		(drawing, 2641, 568, 3900, 800, 0),
		(drawing, 2642, 569, 3900, 800, 0),
		(drawing, 2643, 569, 3900, 800, 0),
		(drawing, 2644, 569, 3900, 800, 0),
		(drawing, 2645, 569, 3900, 800, 0),
		(drawing, 2646, 569, 3900, 800, 0),
		(drawing, 2647, 569, 3900, 800, 0),
		(drawing, 2648, 570, 3900, 800, 0),
		(drawing, 2649, 570, 3900, 800, 0),
		(drawing, 2650, 570, 3900, 800, 0),
		(drawing, 2651, 570, 3900, 800, 0),
		(drawing, 2652, 570, 3900, 800, 0),
		(drawing, 2653, 571, 3900, 800, 0),
		(drawing, 2654, 571, 3900, 800, 0),
		(drawing, 2655, 571, 3900, 800, 0),
		(drawing, 2656, 571, 3900, 800, 0),
		(drawing, 2657, 571, 3900, 800, 0),
		(drawing, 2658, 572, 3900, 800, 0),
		(drawing, 2659, 572, 3900, 800, 0),
		(drawing, 2660, 572, 3900, 800, 0),
		(drawing, 2661, 572, 3900, 800, 0),
		(drawing, 2662, 572, 3900, 800, 0),
		(drawing, 2663, 572, 3900, 800, 0),
		(drawing, 2664, 573, 3900, 800, 0),
		(drawing, 2665, 573, 3900, 800, 0),
		(drawing, 2666, 573, 3900, 800, 0),
		(drawing, 2667, 573, 3900, 800, 0),
		(drawing, 2668, 573, 3900, 800, 0),
		(drawing, 2669, 574, 3900, 800, 0),
		(drawing, 2670, 574, 3900, 800, 0),
		(drawing, 2671, 574, 3900, 800, 0),
		(drawing, 2672, 574, 3900, 800, 0),
		(drawing, 2673, 574, 3900, 800, 0),
		(drawing, 2674, 574, 3900, 800, 0),
		(drawing, 2675, 575, 3900, 800, 0),
		(drawing, 2676, 575, 3900, 800, 0),
		(drawing, 2677, 575, 3900, 800, 0),
		(drawing, 2678, 575, 3900, 800, 0),
		(drawing, 2679, 575, 3900, 800, 0),
		(drawing, 2680, 576, 3900, 800, 0),
		(drawing, 2681, 576, 3900, 800, 0),
		(drawing, 2682, 576, 3900, 800, 0),
		(drawing, 2683, 576, 3900, 800, 0),
		(drawing, 2684, 576, 3900, 800, 0),
		(drawing, 2685, 576, 3900, 800, 0),
		(drawing, 2686, 577, 3900, 800, 0),
		(drawing, 2687, 577, 3900, 800, 0),
		(drawing, 2688, 577, 3900, 800, 0),
		(drawing, 2689, 577, 3900, 800, 0),
		(drawing, 2690, 577, 3900, 800, 0),
		(drawing, 2691, 578, 3900, 800, 0),
		(drawing, 2692, 578, 3900, 800, 0),
		(drawing, 2693, 578, 3900, 800, 0),
		(drawing, 2694, 578, 3900, 800, 0),
		(drawing, 2695, 578, 3900, 800, 0),
		(drawing, 2696, 579, 3900, 800, 0),
		(drawing, 2697, 579, 3900, 800, 0),
		(drawing, 2698, 579, 3900, 800, 0),
		(drawing, 2699, 579, 3900, 800, 0),
		(drawing, 2700, 579, 3900, 800, 0),
		(drawing, 2701, 579, 3900, 800, 0),
		(drawing, 2702, 580, 3900, 800, 0),
		(drawing, 2703, 580, 3900, 800, 0),
		(drawing, 2704, 580, 3900, 800, 0),
		(drawing, 2705, 580, 3900, 800, 0),
		(drawing, 2706, 580, 3900, 800, 0),
		(drawing, 2707, 581, 3900, 800, 0),
		(drawing, 2708, 581, 3900, 800, 0),
		(drawing, 2709, 581, 3900, 800, 0),
		(drawing, 2710, 581, 3900, 800, 0),
		(drawing, 2711, 581, 3900, 800, 0),
		(drawing, 2712, 581, 3900, 800, 0),
		(drawing, 2713, 582, 3900, 800, 0),
		(drawing, 2714, 582, 3900, 800, 0),
		(drawing, 2715, 582, 3900, 800, 0),
		(drawing, 2716, 582, 3900, 800, 0),
		(drawing, 2717, 582, 3900, 800, 0),
		(drawing, 2718, 583, 3900, 800, 0),
		(drawing, 2719, 583, 3900, 800, 0),
		(drawing, 2720, 583, 3900, 800, 0),
		(drawing, 2721, 583, 3900, 800, 0),
		(drawing, 2722, 583, 3900, 800, 0),
		(drawing, 2723, 583, 3900, 800, 0),
		(drawing, 2724, 584, 3900, 800, 0),
		(drawing, 2725, 584, 3900, 800, 0),
		(drawing, 2726, 584, 3900, 800, 0),
		(drawing, 2727, 584, 3900, 800, 0),
		(drawing, 2728, 584, 3900, 800, 0),
		(drawing, 2729, 585, 3900, 800, 0),
		(drawing, 2730, 585, 3900, 800, 0),
		(drawing, 2731, 585, 3900, 800, 0),
		(drawing, 2732, 585, 3900, 800, 0),
		(drawing, 2733, 585, 3900, 800, 0),
		(drawing, 2734, 586, 3900, 800, 0),
		(drawing, 2735, 586, 3900, 800, 0),
		(drawing, 2736, 586, 3900, 800, 0),
		(drawing, 2737, 586, 3900, 800, 0),
		(drawing, 2738, 586, 3900, 800, 0),
		(drawing, 2739, 586, 3900, 800, 0),
		(drawing, 2740, 587, 3900, 800, 0),
		(drawing, 2741, 587, 3900, 800, 0),
		(drawing, 2742, 587, 3900, 800, 0),
		(drawing, 2743, 587, 3900, 800, 0),
		(drawing, 2744, 587, 3900, 800, 0),
		(drawing, 2745, 588, 3900, 800, 0),
		(drawing, 2746, 588, 3900, 800, 0),
		(drawing, 2747, 588, 3900, 800, 0),
		(drawing, 2748, 588, 3900, 800, 0),
		(drawing, 2749, 588, 3900, 800, 0),
		(drawing, 2750, 588, 3900, 800, 0),
		(drawing, 2751, 589, 3900, 800, 0),
		(drawing, 2752, 589, 3900, 800, 0),
		(drawing, 2753, 589, 3900, 800, 0),
		(drawing, 2754, 589, 3900, 800, 0),
		(drawing, 2755, 589, 3900, 800, 0),
		(drawing, 2756, 590, 3900, 800, 0),
		(drawing, 2757, 590, 3900, 800, 0),
		(drawing, 2758, 590, 3900, 800, 0),
		(drawing, 2759, 590, 3900, 800, 0),
		(drawing, 2760, 590, 3900, 800, 0),
		(drawing, 2761, 590, 3900, 800, 0),
		(drawing, 2762, 591, 3900, 800, 0),
		(drawing, 2763, 591, 3900, 800, 0),
		(drawing, 2764, 591, 3900, 800, 0),
		(drawing, 2765, 591, 3900, 800, 0),
		(drawing, 2766, 591, 3900, 800, 0),
		(drawing, 2767, 592, 3900, 800, 0),
		(drawing, 2768, 592, 3900, 800, 0),
		(drawing, 2769, 592, 3900, 800, 0),
		(drawing, 2770, 592, 3900, 800, 0),
		(drawing, 2771, 592, 3900, 800, 0),
		(drawing, 2772, 592, 3900, 800, 0),
		(drawing, 2773, 593, 3900, 800, 0),
		(drawing, 2774, 593, 3900, 800, 0),
		(drawing, 2775, 593, 3900, 800, 0),
		(drawing, 2776, 593, 3900, 800, 0),
		(drawing, 2777, 593, 3900, 800, 0),
		(drawing, 2778, 594, 3900, 800, 0),
		(drawing, 2779, 594, 3900, 800, 0),
		(drawing, 2780, 594, 3900, 800, 0),
		(drawing, 2781, 594, 3900, 800, 0),
		(drawing, 2782, 594, 3900, 800, 0),
		(drawing, 2783, 595, 3900, 800, 0),
		(drawing, 2784, 595, 3900, 800, 0),
		(drawing, 2785, 595, 3900, 800, 0),
		(drawing, 2786, 595, 3900, 800, 0),
		(drawing, 2787, 595, 3900, 800, 0),
		(drawing, 2788, 595, 3900, 800, 0),
		(drawing, 2789, 596, 3900, 800, 0),
		(drawing, 2790, 596, 3900, 800, 0),
		(drawing, 2791, 596, 3900, 800, 0),
		(drawing, 2792, 596, 3900, 800, 0),
		(drawing, 2793, 596, 3900, 800, 0),
		(drawing, 2794, 597, 3900, 800, 0),
		(drawing, 2795, 597, 3900, 800, 0),
		(drawing, 2796, 597, 3900, 800, 0),
		(drawing, 2797, 597, 3900, 800, 0),
		(drawing, 2798, 597, 3900, 800, 0),
		(drawing, 2799, 597, 3900, 800, 0),
		(drawing, 2800, 598, 3900, 800, 0),
		(drawing, 2801, 598, 3900, 800, 0),
		(drawing, 2802, 598, 3900, 800, 0),
		(drawing, 2803, 598, 3900, 800, 0),
		(drawing, 2804, 598, 3900, 800, 0),
		(drawing, 2805, 599, 3900, 800, 0),
		(drawing, 2806, 599, 3900, 800, 0),
		(drawing, 2807, 599, 3900, 800, 0),
		(drawing, 2808, 599, 3900, 800, 0),
		(drawing, 2809, 599, 3900, 800, 0),
		(drawing, 2810, 599, 3900, 800, 0),
		(drawing, 2811, 600, 3900, 800, 0),
		(drawing, 2812, 600, 3900, 800, 0),
		(drawing, 2813, 600, 3900, 800, 0),
		(drawing, 2814, 600, 3900, 800, 0),
		(drawing, 2815, 600, 3900, 800, 0),
		(drawing, 2816, 601, 3900, 800, 0),
		(drawing, 2817, 601, 3900, 800, 0),
		(drawing, 2818, 601, 3900, 800, 0),
		(drawing, 2819, 601, 3900, 800, 0),
		(drawing, 2820, 601, 3900, 800, 0),
		(drawing, 2821, 602, 3900, 800, 0),
		(drawing, 2822, 602, 3900, 800, 0),
		(drawing, 2823, 602, 3900, 800, 0),
		(drawing, 2824, 602, 3900, 800, 0),
		(drawing, 2825, 602, 3900, 800, 0),
		(drawing, 2826, 602, 3900, 800, 0),
		(drawing, 2827, 603, 3900, 800, 0),
		(drawing, 2828, 603, 3900, 800, 0),
		(drawing, 2829, 603, 3900, 800, 0),
		(drawing, 2830, 603, 3900, 800, 0),
		(drawing, 2831, 603, 3900, 800, 0),
		(drawing, 2832, 604, 3900, 800, 0),
		(drawing, 2833, 604, 3900, 800, 0),
		(drawing, 2834, 604, 3900, 800, 0),
		(drawing, 2835, 604, 3900, 800, 0),
		(drawing, 2836, 604, 3900, 800, 0),
		(drawing, 2837, 604, 3900, 800, 0),
		(drawing, 2838, 605, 3900, 800, 0),
		(drawing, 2839, 605, 3900, 800, 0),
		(drawing, 2840, 605, 3900, 800, 0),
		(drawing, 2841, 605, 3900, 800, 0),
		(drawing, 2842, 605, 3900, 800, 0),
		(drawing, 2843, 606, 3900, 800, 0),
		(drawing, 2844, 606, 3900, 800, 0),
		(drawing, 2845, 606, 3900, 800, 0),
		(drawing, 2846, 606, 3900, 800, 0),
		(drawing, 2847, 606, 3900, 800, 0),
		(drawing, 2848, 606, 3900, 800, 0),
		(drawing, 2849, 607, 3900, 800, 0),
		(drawing, 2850, 607, 3900, 800, 0),
		(drawing, 2851, 607, 3900, 800, 0),
		(drawing, 2852, 607, 3900, 800, 0),
		(drawing, 2853, 607, 3900, 800, 0),
		(drawing, 2854, 608, 3900, 800, 0),
		(drawing, 2855, 608, 3900, 800, 0),
		(drawing, 2856, 608, 3900, 800, 0),
		(drawing, 2857, 608, 3900, 800, 0),
		(drawing, 2858, 608, 3900, 800, 0),
		(drawing, 2859, 608, 3900, 800, 0),
		(drawing, 2860, 609, 3900, 800, 0),
		(drawing, 2861, 609, 3900, 800, 0),
		(drawing, 2862, 609, 3900, 800, 0),
		(drawing, 2863, 609, 3900, 800, 0),
		(drawing, 2864, 609, 3900, 800, 0),
		(drawing, 2865, 610, 3900, 800, 0),
		(drawing, 2866, 610, 3900, 800, 0),
		(drawing, 2867, 610, 3900, 800, 0),
		(drawing, 2868, 610, 3900, 800, 0),
		(drawing, 2869, 610, 3900, 800, 0),
		(drawing, 2870, 611, 3900, 800, 0),
		(drawing, 2871, 611, 3900, 800, 0),
		(drawing, 2872, 611, 3900, 800, 0),
		(drawing, 2873, 611, 3900, 800, 0),
		(drawing, 2874, 611, 3900, 800, 0),
		(drawing, 2875, 611, 3900, 800, 0),
		(drawing, 2876, 612, 3900, 800, 0),
		(drawing, 2877, 612, 3900, 800, 0),
		(drawing, 2878, 612, 3900, 800, 0),
		(drawing, 2879, 612, 3900, 800, 0),
		(drawing, 2880, 612, 3900, 800, 0),
		(drawing, 2881, 613, 3900, 800, 0),
		(drawing, 2882, 613, 3900, 800, 0),
		(drawing, 2883, 613, 3900, 800, 0),
		(drawing, 2884, 613, 3900, 800, 0),
		(drawing, 2885, 613, 3900, 800, 0),
		(drawing, 2886, 613, 3900, 800, 0),
		(drawing, 2887, 614, 3900, 800, 0),
		(drawing, 2888, 614, 3900, 800, 0),
		(drawing, 2889, 614, 3900, 800, 0),
		(drawing, 2890, 614, 3900, 800, 0),
		(drawing, 2891, 614, 3900, 800, 0),
		(drawing, 2892, 615, 3900, 800, 0),
		(drawing, 2893, 615, 3900, 800, 0),
		(drawing, 2894, 615, 3900, 800, 0),
		(drawing, 2895, 615, 3900, 800, 0),
		(drawing, 2896, 615, 3900, 800, 0),
		(drawing, 2897, 615, 3900, 800, 0),
		(drawing, 2898, 616, 3900, 800, 0),
		(drawing, 2899, 616, 3900, 800, 0),
		(drawing, 2900, 616, 3900, 800, 0),
		(drawing, 2901, 616, 3900, 800, 0),
		(drawing, 2902, 616, 3900, 800, 0),
		(drawing, 2903, 617, 3900, 800, 0),
		(drawing, 2904, 617, 3900, 800, 0),
		(drawing, 2905, 617, 3900, 800, 0),
		(drawing, 2906, 617, 3900, 800, 0),
		(drawing, 2907, 617, 3900, 800, 0),
		(drawing, 2908, 618, 3900, 800, 0),
		(drawing, 2909, 618, 3900, 800, 0),
		(drawing, 2910, 618, 3900, 800, 0),
		(drawing, 2911, 618, 3900, 800, 0),
		(drawing, 2912, 618, 3900, 800, 0),
		(drawing, 2913, 618, 3900, 800, 0),
		(drawing, 2914, 619, 3900, 800, 0),
		(drawing, 2915, 619, 3900, 800, 0),
		(drawing, 2916, 619, 3900, 800, 0),
		(drawing, 2917, 619, 3900, 800, 0),
		(drawing, 2918, 619, 3900, 800, 0),
		(drawing, 2919, 620, 3900, 800, 0),
		(drawing, 2920, 620, 3900, 800, 0),
		(drawing, 2921, 620, 3900, 800, 0),
		(drawing, 2922, 620, 3900, 800, 0),
		(drawing, 2923, 620, 3900, 800, 0),
		(drawing, 2924, 620, 3900, 800, 0),
		(drawing, 2925, 621, 3900, 800, 0),
		(drawing, 2926, 621, 3900, 800, 0),
		(drawing, 2927, 621, 3900, 800, 0),
		(drawing, 2928, 621, 3900, 800, 0),
		(drawing, 2929, 621, 3900, 800, 0),
		(drawing, 2930, 622, 3900, 800, 0),
		(drawing, 2931, 622, 3900, 800, 0),
		(drawing, 2932, 622, 3900, 800, 0),
		(drawing, 2933, 622, 3900, 800, 0),
		(drawing, 2934, 622, 3900, 800, 0),
		(drawing, 2935, 622, 3900, 800, 0),
		(drawing, 2936, 623, 3900, 800, 0),
		(drawing, 2937, 623, 3900, 800, 0),
		(drawing, 2938, 623, 3900, 800, 0),
		(drawing, 2939, 623, 3900, 800, 0),
		(drawing, 2940, 623, 3900, 800, 0),
		(drawing, 2941, 624, 3900, 800, 0),
		(drawing, 2942, 624, 3900, 800, 0),
		(drawing, 2943, 624, 3900, 800, 0),
		(drawing, 2944, 624, 3900, 800, 0),
		(drawing, 2945, 624, 3900, 800, 0),
		(drawing, 2946, 625, 3900, 800, 0),
		(drawing, 2947, 625, 3900, 800, 0),
		(drawing, 2948, 625, 3900, 800, 0),
		(drawing, 2949, 625, 3900, 800, 0),
		(drawing, 2950, 625, 3900, 800, 0),
		(drawing, 2951, 625, 3900, 800, 0),
		(drawing, 2952, 626, 3900, 800, 0),
		(drawing, 2953, 626, 3900, 800, 0),
		(drawing, 2954, 626, 3900, 800, 0),
		(drawing, 2955, 626, 3900, 800, 0),
		(drawing, 2956, 626, 3900, 800, 0),
		(drawing, 2957, 627, 3900, 800, 0),
		(drawing, 2958, 627, 3900, 800, 0),
		(drawing, 2959, 627, 3900, 800, 0),
		(drawing, 2960, 627, 3900, 800, 0),
		(drawing, 2961, 627, 3900, 800, 0),
		(drawing, 2962, 627, 3900, 800, 0),
		(drawing, 2963, 628, 3900, 800, 0),
		(drawing, 2964, 628, 3900, 800, 0),
		(drawing, 2965, 628, 3900, 800, 0),
		(drawing, 2966, 628, 3900, 800, 0),
		(drawing, 2967, 628, 3900, 800, 0),
		(drawing, 2968, 629, 3900, 800, 0),
		(drawing, 2969, 629, 3900, 800, 0),
		(drawing, 2970, 629, 3900, 800, 0),
		(drawing, 2971, 629, 3900, 800, 0),
		(drawing, 2972, 629, 3900, 800, 0),
		(drawing, 2973, 629, 3900, 800, 0),
		(drawing, 2974, 630, 3900, 800, 0),
		(drawing, 2975, 630, 3900, 800, 0),
		(drawing, 2976, 630, 3900, 800, 0),
		(drawing, 2977, 630, 3900, 800, 0),
		(drawing, 2978, 630, 3900, 800, 0),
		(drawing, 2979, 631, 3900, 800, 0),
		(drawing, 2980, 631, 3900, 800, 0),
		(drawing, 2981, 631, 3900, 800, 0),
		(drawing, 2982, 631, 3900, 800, 0),
		(drawing, 2983, 631, 3900, 800, 0),
		(drawing, 2984, 631, 3900, 800, 0),
		(drawing, 2985, 632, 3900, 800, 0),
		(drawing, 2986, 632, 3900, 800, 0),
		(drawing, 2987, 632, 3900, 800, 0),
		(drawing, 2988, 632, 3900, 800, 0),
		(drawing, 2989, 632, 3900, 800, 0),
		(drawing, 2990, 633, 3900, 800, 0),
		(drawing, 2991, 633, 3900, 800, 0),
		(drawing, 2992, 633, 3900, 800, 0),
		(drawing, 2993, 633, 3900, 800, 0),
		(drawing, 2994, 633, 3900, 800, 0),
		(drawing, 2995, 634, 3900, 800, 0),
		(drawing, 2996, 634, 3900, 800, 0),
		(drawing, 2997, 634, 3900, 800, 0),
		(drawing, 2998, 634, 3900, 800, 0),
		(drawing, 2999, 634, 3900, 800, 0),
		(drawing, 3000, 634, 3900, 800, 0),
		(drawing, 3001, 635, 3900, 800, 0),
		(drawing, 3002, 635, 3900, 800, 0),
		(drawing, 3003, 635, 3900, 800, 0),
		(drawing, 3004, 635, 3900, 800, 0),
		(drawing, 3005, 635, 3900, 800, 0),
		(drawing, 3006, 636, 3900, 800, 0),
		(drawing, 3007, 636, 3900, 800, 0),
		(drawing, 3008, 636, 3900, 800, 0),
		(drawing, 3009, 636, 3900, 800, 0),
		(drawing, 3010, 636, 3900, 800, 0),
		(drawing, 3011, 636, 3900, 800, 0),
		(drawing, 3012, 637, 3900, 800, 0),
		(drawing, 3013, 637, 3900, 800, 0),
		(drawing, 3014, 637, 3900, 800, 0),
		(drawing, 3015, 637, 3900, 800, 0),
		(drawing, 3016, 637, 3900, 800, 0),
		(drawing, 3017, 638, 3900, 800, 0),
		(drawing, 3018, 638, 3900, 800, 0),
		(drawing, 3019, 638, 3900, 800, 0),
		(drawing, 3020, 638, 3900, 800, 0),
		(drawing, 3021, 638, 3900, 800, 0),
		(drawing, 3022, 638, 3900, 800, 0),
		(drawing, 3023, 639, 3900, 800, 0),
		(drawing, 3024, 639, 3900, 800, 0),
		(drawing, 3025, 639, 3900, 800, 0),
		(drawing, 3026, 639, 3900, 800, 0),
		(drawing, 3027, 639, 3900, 800, 0),
		(drawing, 3028, 640, 3900, 800, 0),
		(drawing, 3029, 640, 3900, 800, 0),
		(drawing, 3030, 640, 3900, 800, 0),
		(drawing, 3031, 640, 3900, 800, 0),
		(drawing, 3032, 640, 3900, 800, 0),
		(drawing, 3033, 641, 3900, 800, 0),
		(drawing, 3034, 641, 3900, 800, 0),
		(drawing, 3035, 641, 3900, 800, 0),
		(drawing, 3036, 641, 3900, 800, 0),
		(drawing, 3037, 641, 3900, 800, 0),
		(drawing, 3038, 641, 3900, 800, 0),
		(drawing, 3039, 642, 3900, 800, 0),
		(drawing, 3040, 642, 3900, 800, 0),
		(drawing, 3041, 642, 3900, 800, 0),
		(drawing, 3042, 642, 3900, 800, 0),
		(drawing, 3043, 642, 3900, 800, 0),
		(drawing, 3044, 643, 3900, 800, 0),
		(drawing, 3045, 643, 3900, 800, 0),
		(drawing, 3046, 643, 3900, 800, 0),
		(drawing, 3047, 643, 3900, 800, 0),
		(drawing, 3048, 643, 3900, 800, 0),
		(drawing, 3049, 643, 3900, 800, 0),
		(drawing, 3050, 644, 3900, 800, 0),
		(drawing, 3051, 644, 3900, 800, 0),
		(drawing, 3052, 644, 3900, 800, 0),
		(drawing, 3053, 644, 3900, 800, 0),
		(drawing, 3054, 644, 3900, 800, 0),
		(drawing, 3055, 645, 3900, 800, 0),
		(drawing, 3056, 645, 3900, 800, 0),
		(drawing, 3057, 645, 3900, 800, 0),
		(drawing, 3058, 645, 3900, 800, 0),
		(drawing, 3059, 645, 3900, 800, 0),
		(drawing, 3060, 645, 3900, 800, 0),
		(drawing, 3061, 646, 3900, 800, 0),
		(drawing, 3062, 646, 3900, 800, 0),
		(drawing, 3063, 646, 3900, 800, 0),
		(drawing, 3064, 646, 3900, 800, 0),
		(drawing, 3065, 646, 3900, 800, 0),
		(drawing, 3066, 647, 3900, 800, 0),
		(drawing, 3067, 647, 3900, 800, 0),
		(drawing, 3068, 647, 3900, 800, 0),
		(drawing, 3069, 647, 3900, 800, 0),
		(drawing, 3070, 647, 3900, 800, 0),
		(drawing, 3071, 647, 3900, 800, 0),
		(drawing, 3072, 648, 3900, 800, 0),
		(drawing, 3073, 648, 3900, 800, 0),
		(drawing, 3074, 648, 3900, 800, 0),
		(drawing, 3075, 648, 3900, 800, 0),
		(drawing, 3076, 648, 3900, 800, 0),
		(drawing, 3077, 649, 3900, 800, 0),
		(drawing, 3078, 649, 3900, 800, 0),
		(drawing, 3079, 649, 3900, 800, 0),
		(drawing, 3080, 649, 3900, 800, 0),
		(drawing, 3081, 649, 3900, 800, 0),
		(drawing, 3082, 650, 3900, 800, 0),
		(drawing, 3083, 650, 3900, 800, 0),
		(drawing, 3084, 650, 3900, 800, 0),
		(drawing, 3085, 650, 3900, 800, 0),
		(drawing, 3086, 650, 3900, 800, 0),
		(drawing, 3087, 650, 3900, 800, 0),
		(drawing, 3088, 651, 3900, 800, 0),
		(drawing, 3089, 651, 3900, 800, 0),
		(drawing, 3090, 651, 3900, 800, 0),
		(drawing, 3091, 651, 3900, 800, 0),
		(drawing, 3092, 651, 3900, 800, 0),
		(drawing, 3093, 652, 3900, 800, 0),
		(drawing, 3094, 652, 3900, 800, 0),
		(drawing, 3095, 652, 3900, 800, 0),
		(drawing, 3096, 652, 3900, 800, 0),
		(drawing, 3097, 652, 3900, 800, 0),
		(drawing, 3098, 652, 3900, 800, 0),
		(drawing, 3099, 653, 3900, 800, 0),
		(drawing, 3100, 653, 3900, 800, 0),
		(drawing, 3101, 653, 3900, 800, 0),
		(drawing, 3102, 653, 3900, 800, 0),
		(drawing, 3103, 653, 3900, 800, 0),
		(drawing, 3104, 654, 3900, 800, 0),
		(drawing, 3105, 654, 3900, 800, 0),
		(drawing, 3106, 654, 3900, 800, 0),
		(drawing, 3107, 654, 3900, 800, 0),
		(drawing, 3108, 654, 3900, 800, 0),
		(drawing, 3109, 654, 3900, 800, 0),
		(drawing, 3110, 655, 3900, 800, 0),
		(drawing, 3111, 655, 3900, 800, 0),
		(drawing, 3112, 655, 3900, 800, 0),
		(drawing, 3113, 655, 3900, 800, 0),
		(drawing, 3114, 655, 3900, 800, 0),
		(drawing, 3115, 656, 3900, 800, 0),
		(drawing, 3116, 656, 3900, 800, 0),
		(drawing, 3117, 656, 3900, 800, 0),
		(drawing, 3118, 656, 3900, 800, 0),
		(drawing, 3119, 656, 3900, 800, 0),
		(drawing, 3120, 657, 3900, 800, 0),
		(drawing, 3121, 657, 3900, 800, 0),
		(drawing, 3122, 657, 3900, 800, 0),
		(drawing, 3123, 657, 3900, 800, 0),
		(drawing, 3124, 657, 3900, 800, 0),
		(drawing, 3125, 657, 3900, 800, 0),
		(drawing, 3126, 658, 3900, 800, 0),
		(drawing, 3127, 658, 3900, 800, 0),
		(drawing, 3128, 658, 3900, 800, 0),
		(drawing, 3129, 658, 3900, 800, 0),
		(drawing, 3130, 658, 3900, 800, 0),
		(drawing, 3131, 659, 3900, 800, 0),
		(drawing, 3132, 659, 3900, 800, 0),
		(drawing, 3133, 659, 3900, 800, 0),
		(drawing, 3134, 659, 3900, 800, 0),
		(drawing, 3135, 659, 3900, 800, 0),
		(drawing, 3136, 659, 3900, 800, 0),
		(drawing, 3137, 660, 3900, 800, 0),
		(drawing, 3138, 660, 3900, 800, 0),
		(drawing, 3139, 660, 3900, 800, 0),
		(drawing, 3140, 660, 3900, 800, 0),
		(drawing, 3141, 660, 3900, 800, 0),
		(drawing, 3142, 661, 3900, 800, 0),
		(drawing, 3143, 661, 3900, 800, 0),
		(drawing, 3144, 661, 3900, 800, 0),
		(drawing, 3145, 661, 3900, 800, 0),
		(drawing, 3146, 661, 3900, 800, 0),
		(drawing, 3147, 661, 3900, 800, 0),
		(drawing, 3148, 662, 3900, 800, 0),
		(drawing, 3149, 662, 3900, 800, 0),
		(drawing, 3150, 662, 3900, 800, 0),
		(drawing, 3151, 662, 3900, 800, 0),
		(drawing, 3152, 662, 3900, 800, 0),
		(drawing, 3153, 663, 3900, 800, 0),
		(drawing, 3154, 663, 3900, 800, 0),
		(drawing, 3155, 663, 3900, 800, 0),
		(drawing, 3156, 663, 3900, 800, 0),
		(drawing, 3157, 663, 3900, 800, 0),
		(drawing, 3158, 664, 3900, 800, 0),
		(drawing, 3159, 664, 3900, 800, 0),
		(drawing, 3160, 664, 3900, 800, 0),
		(drawing, 3161, 664, 3900, 800, 0),
		(drawing, 3162, 664, 3900, 800, 0),
		(drawing, 3163, 664, 3900, 800, 0),
		(drawing, 3164, 665, 3900, 800, 0),
		(drawing, 3165, 665, 3900, 800, 0),
		(drawing, 3166, 665, 3900, 800, 0),
		(drawing, 3167, 665, 3900, 800, 0),
		(drawing, 3168, 665, 3900, 800, 0),
		(drawing, 3169, 666, 3900, 800, 0),
		(drawing, 3170, 666, 3900, 800, 0),
		(drawing, 3171, 666, 3900, 800, 0),
		(drawing, 3172, 666, 3900, 800, 0),
		(drawing, 3173, 666, 3900, 800, 0),
		(drawing, 3174, 666, 3900, 800, 0),
		(drawing, 3175, 667, 3900, 800, 0),
		(drawing, 3176, 667, 3900, 800, 0),
		(drawing, 3177, 667, 3900, 800, 0),
		(drawing, 3178, 667, 3900, 800, 0),
		(drawing, 3179, 667, 3900, 800, 0),
		(drawing, 3180, 668, 3900, 800, 0),
		(drawing, 3181, 668, 3900, 800, 0),
		(drawing, 3182, 668, 3900, 800, 0),
		(drawing, 3183, 668, 3900, 800, 0),
		(drawing, 3184, 668, 3900, 800, 0),
		(drawing, 3185, 668, 3900, 800, 0),
		(drawing, 3186, 669, 3900, 800, 0),
		(drawing, 3187, 669, 3900, 800, 0),
		(drawing, 3188, 669, 3900, 800, 0),
		(drawing, 3189, 669, 3900, 800, 0),
		(drawing, 3190, 669, 3900, 800, 0),
		(drawing, 3191, 670, 3900, 800, 0),
		(drawing, 3192, 670, 3900, 800, 0),
		(drawing, 3193, 670, 3900, 800, 0),
		(drawing, 3194, 670, 3900, 800, 0),
		(drawing, 3195, 670, 3900, 800, 0),
		(drawing, 3196, 670, 3900, 800, 0),
		(drawing, 3197, 671, 3900, 800, 0),
		(drawing, 3198, 671, 3900, 800, 0),
		(drawing, 3199, 671, 3900, 800, 0),
		(drawing, 3200, 671, 3900, 800, 0),
		(drawing, 3201, 671, 3900, 800, 0),
		(drawing, 3202, 672, 3900, 800, 0),
		(drawing, 3203, 672, 3900, 800, 0),
		(drawing, 3204, 672, 3900, 800, 0),
		(drawing, 3205, 672, 3900, 800, 0),
		(drawing, 3206, 672, 3900, 800, 0),
		(drawing, 3207, 673, 3900, 800, 0),
		(drawing, 3208, 673, 3900, 800, 0),
		(drawing, 3209, 673, 3900, 800, 0),
		(drawing, 3210, 673, 3900, 800, 0),
		(drawing, 3211, 673, 3900, 800, 0),
		(drawing, 3212, 673, 3900, 800, 0),
		(drawing, 3213, 674, 3900, 800, 0),
		(drawing, 3214, 674, 3900, 800, 0),
		(drawing, 3215, 674, 3900, 800, 0),
		(drawing, 3216, 674, 3900, 800, 0),
		(drawing, 3217, 674, 3900, 800, 0),
		(drawing, 3218, 675, 3900, 800, 0),
		(drawing, 3219, 675, 3900, 800, 0),
		(drawing, 3220, 675, 3900, 800, 0),
		(drawing, 3221, 675, 3900, 800, 0),
		(drawing, 3222, 675, 3900, 800, 0),
		(drawing, 3223, 675, 3900, 800, 0),
		(drawing, 3224, 676, 3900, 800, 0),
		(drawing, 3225, 676, 3900, 800, 0),
		(drawing, 3226, 676, 3900, 800, 0),
		(drawing, 3227, 676, 3900, 800, 0),
		(drawing, 3228, 676, 3900, 800, 0),
		(drawing, 3229, 677, 3900, 800, 0),
		(drawing, 3230, 677, 3900, 800, 0),
		(drawing, 3231, 677, 3900, 800, 0),
		(drawing, 3232, 677, 3900, 800, 0),
		(drawing, 3233, 677, 3900, 800, 0),
		(drawing, 3234, 677, 3900, 800, 0),
		(drawing, 3235, 678, 3900, 800, 0),
		(drawing, 3236, 678, 3900, 800, 0),
		(drawing, 3237, 678, 3900, 800, 0),
		(drawing, 3238, 678, 3900, 800, 0),
		(drawing, 3239, 678, 3900, 800, 0),
		(drawing, 3240, 679, 3900, 800, 0),
		(drawing, 3241, 679, 3900, 800, 0),
		(drawing, 3242, 679, 3900, 800, 0),
		(drawing, 3243, 679, 3900, 800, 0),
		(drawing, 3244, 679, 3900, 800, 0),
		(drawing, 3245, 680, 3900, 800, 0),
		(drawing, 3246, 680, 3900, 800, 0),
		(drawing, 3247, 680, 3900, 800, 0),
		(drawing, 3248, 680, 3900, 800, 0),
		(drawing, 3249, 680, 3900, 800, 0),
		(drawing, 3250, 680, 3900, 800, 0),
		(drawing, 3251, 681, 3900, 800, 0),
		(drawing, 3252, 681, 3900, 800, 0),
		(drawing, 3253, 681, 3900, 800, 0),
		(drawing, 3254, 681, 3900, 800, 0),
		(drawing, 3255, 681, 3900, 800, 0),
		(drawing, 3256, 682, 3900, 800, 0),
		(drawing, 3257, 682, 3900, 800, 0),
		(drawing, 3258, 682, 3900, 800, 0),
		(drawing, 3259, 682, 3900, 800, 0),
		(drawing, 3260, 682, 3900, 800, 0),
		(drawing, 3261, 682, 3900, 800, 0),
		(drawing, 3262, 683, 3900, 800, 0),
		(drawing, 3263, 683, 3900, 800, 0),
		(drawing, 3264, 683, 3900, 800, 0),
		(drawing, 3265, 683, 3900, 800, 0),
		(drawing, 3266, 683, 3900, 800, 0),
		(drawing, 3267, 684, 3900, 800, 0),
		(drawing, 3268, 684, 3900, 800, 0),
		(drawing, 3269, 684, 3900, 800, 0),
		(drawing, 3270, 684, 3900, 800, 0),
		(drawing, 3271, 684, 3900, 800, 0),
		(drawing, 3272, 684, 3900, 800, 0),
		(drawing, 3273, 685, 3900, 800, 0),
		(drawing, 3274, 685, 3900, 800, 0),
		(drawing, 3275, 685, 3900, 800, 0),
		(drawing, 3276, 685, 3900, 800, 0),
		(drawing, 3277, 685, 3900, 800, 0),
		(drawing, 3278, 686, 3900, 800, 0),
		(drawing, 3279, 686, 3900, 800, 0),
		(drawing, 3280, 686, 3900, 800, 0),
		(drawing, 3281, 686, 3900, 800, 0),
		(drawing, 3282, 686, 3900, 800, 0),
		(drawing, 3283, 686, 3900, 800, 0),
		(drawing, 3284, 687, 3900, 800, 0),
		(drawing, 3285, 687, 3900, 800, 0),
		(drawing, 3286, 687, 3900, 800, 0),
		(drawing, 3287, 687, 3900, 800, 0),
		(drawing, 3288, 687, 3900, 800, 0),
		(drawing, 3289, 688, 3900, 800, 0),
		(drawing, 3290, 688, 3900, 800, 0),
		(drawing, 3291, 688, 3900, 800, 0),
		(drawing, 3292, 688, 3900, 800, 0),
		(drawing, 3293, 688, 3900, 800, 0),
		(drawing, 3294, 689, 3900, 800, 0),
		(drawing, 3295, 689, 3900, 800, 0),
		(drawing, 3296, 689, 3900, 800, 0),
		(drawing, 3297, 689, 3900, 800, 0),
		(drawing, 3298, 689, 3900, 800, 0),
		(drawing, 3299, 689, 3900, 800, 0),
		(drawing, 3300, 690, 3900, 800, 0),
		(drawing, 3301, 690, 3900, 800, 0),
		(drawing, 3302, 690, 3900, 800, 0),
		(drawing, 3303, 690, 3900, 800, 0),
		(drawing, 3304, 690, 3900, 800, 0),
		(drawing, 3305, 691, 3900, 800, 0),
		(drawing, 3306, 691, 3900, 800, 0),
		(drawing, 3307, 691, 3900, 800, 0),
		(drawing, 3308, 691, 3900, 800, 0),
		(drawing, 3309, 691, 3900, 800, 0),
		(drawing, 3310, 691, 3900, 800, 0),
		(drawing, 3311, 692, 3900, 800, 0),
		(drawing, 3312, 692, 3900, 800, 0),
		(drawing, 3313, 692, 3900, 800, 0),
		(drawing, 3314, 692, 3900, 800, 0),
		(drawing, 3315, 692, 3900, 800, 0),
		(drawing, 3316, 693, 3900, 800, 0),
		(drawing, 3317, 693, 3900, 800, 0),
		(drawing, 3318, 693, 3900, 800, 0),
		(drawing, 3319, 693, 3900, 800, 0),
		(drawing, 3320, 693, 3900, 800, 0),
		(drawing, 3321, 693, 3900, 800, 0),
		(drawing, 3322, 694, 3900, 800, 0),
		(drawing, 3323, 694, 3900, 800, 0),
		(drawing, 3324, 694, 3900, 800, 0),
		(drawing, 3325, 694, 3900, 800, 0),
		(drawing, 3326, 694, 3900, 800, 0),
		(drawing, 3327, 695, 3900, 800, 0),
		(drawing, 3328, 695, 3900, 800, 0),
		(drawing, 3329, 695, 3900, 800, 0),
		(drawing, 3330, 695, 3900, 800, 0),
		(drawing, 3331, 695, 3900, 800, 0),
		(drawing, 3332, 696, 3900, 800, 0),
		(drawing, 3333, 696, 3900, 800, 0),
		(drawing, 3334, 696, 3900, 800, 0),
		(drawing, 3335, 696, 3900, 800, 0),
		(drawing, 3336, 696, 3900, 800, 0),
		(drawing, 3337, 696, 3900, 800, 0),
		(drawing, 3338, 697, 3900, 800, 0),
		(drawing, 3339, 697, 3900, 800, 0),
		(drawing, 3340, 697, 3900, 800, 0),
		(drawing, 3341, 697, 3900, 800, 0),
		(drawing, 3342, 697, 3900, 800, 0),
		(drawing, 3343, 698, 3900, 800, 0),
		(drawing, 3344, 698, 3900, 800, 0),
		(drawing, 3345, 698, 3900, 800, 0),
		(drawing, 3346, 698, 3900, 800, 0),
		(drawing, 3347, 698, 3900, 800, 0),
		(drawing, 3348, 698, 3900, 800, 0),
		(drawing, 3349, 699, 3900, 800, 0),
		(drawing, 3350, 699, 3900, 800, 0),
		(drawing, 3351, 699, 3900, 800, 0),
		(drawing, 3352, 699, 3900, 800, 0),
		(drawing, 3353, 699, 3900, 800, 0),
		(drawing, 3354, 700, 3900, 800, 0),
		(drawing, 3355, 700, 3900, 800, 0),
		(drawing, 3356, 700, 3900, 800, 0),
		(drawing, 3357, 700, 3900, 800, 0),
		(drawing, 3358, 700, 3900, 800, 0),
		(drawing, 3359, 700, 3900, 800, 0),
		(drawing, 3360, 701, 3900, 800, 0),
		(drawing, 3361, 701, 3900, 800, 0),
		(drawing, 3362, 701, 3900, 800, 0),
		(drawing, 3363, 701, 3900, 800, 0),
		(drawing, 3364, 701, 3900, 800, 0),
		(drawing, 3365, 702, 3900, 800, 0),
		(drawing, 3366, 702, 3900, 800, 0),
		(drawing, 3367, 702, 3900, 800, 0),
		(drawing, 3368, 702, 3900, 800, 0),
		(drawing, 3369, 702, 3900, 800, 0),
		(drawing, 3370, 703, 3900, 800, 0),
		(drawing, 3371, 703, 3900, 800, 0),
		(drawing, 3372, 703, 3900, 800, 0),
		(drawing, 3373, 703, 3900, 800, 0),
		(drawing, 3374, 703, 3900, 800, 0),
		(drawing, 3375, 703, 3900, 800, 0),
		(drawing, 3376, 704, 3900, 800, 0),
		(drawing, 3377, 704, 3900, 800, 0),
		(drawing, 3378, 704, 3900, 800, 0),
		(drawing, 3379, 704, 3900, 800, 0),
		(drawing, 3380, 704, 3900, 800, 0),
		(drawing, 3381, 705, 3900, 800, 0),
		(drawing, 3382, 705, 3900, 800, 0),
		(drawing, 3383, 705, 3900, 800, 0),
		(drawing, 3384, 705, 3900, 800, 0),
		(drawing, 3385, 705, 3900, 800, 0),
		(drawing, 3386, 705, 3900, 800, 0),
		(drawing, 3387, 706, 3900, 800, 0),
		(drawing, 3388, 706, 3900, 800, 0),
		(drawing, 3389, 706, 3900, 800, 0),
		(drawing, 3390, 706, 3900, 800, 0),
		(drawing, 3391, 706, 3900, 800, 0),
		(drawing, 3392, 707, 3900, 800, 0),
		(drawing, 3393, 707, 3900, 800, 0),
		(drawing, 3394, 707, 3900, 800, 0),
		(drawing, 3395, 707, 3900, 800, 0),
		(drawing, 3396, 707, 3900, 800, 0),
		(drawing, 3397, 707, 3900, 800, 0),
		(drawing, 3398, 708, 3900, 800, 0),
		(drawing, 3399, 708, 3900, 800, 0),
		(drawing, 3400, 708, 3900, 800, 0),
		(drawing, 3401, 708, 3900, 800, 0),
		(drawing, 3402, 708, 3900, 800, 0),
		(drawing, 3403, 709, 3900, 800, 0),
		(drawing, 3404, 709, 3900, 800, 0),
		(drawing, 3405, 709, 3900, 800, 0),
		(drawing, 3406, 709, 3900, 800, 0),
		(drawing, 3407, 709, 3900, 800, 0),
		(drawing, 3408, 709, 3900, 800, 0),
		(drawing, 3409, 710, 3900, 800, 0),
		(drawing, 3410, 710, 3900, 800, 0),
		(drawing, 3411, 710, 3900, 800, 0),
		(drawing, 3412, 710, 3900, 800, 0),
		(drawing, 3413, 710, 3900, 800, 0),
		(drawing, 3414, 711, 3900, 800, 0),
		(drawing, 3415, 711, 3900, 800, 0),
		(drawing, 3416, 711, 3900, 800, 0),
		(drawing, 3417, 711, 3900, 800, 0),
		(drawing, 3418, 711, 3900, 800, 0),
		(drawing, 3419, 712, 3900, 800, 0),
		(drawing, 3420, 712, 3900, 800, 0),
		(drawing, 3421, 712, 3900, 800, 0),
		(drawing, 3422, 712, 3900, 800, 0),
		(drawing, 3423, 712, 3900, 800, 0),
		(drawing, 3424, 712, 3900, 800, 0),
		(drawing, 3425, 713, 3900, 800, 0),
		(drawing, 3426, 713, 3900, 800, 0),
		(drawing, 3427, 713, 3900, 800, 0),
		(drawing, 3428, 713, 3900, 800, 0),
		(drawing, 3429, 713, 3900, 800, 0),
		(drawing, 3430, 714, 3900, 800, 0),
		(drawing, 3431, 714, 3900, 800, 0),
		(drawing, 3432, 714, 3900, 800, 0),
		(drawing, 3433, 714, 3900, 800, 0),
		(drawing, 3434, 714, 3900, 800, 0),
		(drawing, 3435, 714, 3900, 800, 0),
		(drawing, 3436, 715, 3900, 800, 0),
		(drawing, 3437, 715, 3900, 800, 0),
		(drawing, 3438, 715, 3900, 800, 0),
		(drawing, 3439, 715, 3900, 800, 0),
		(drawing, 3440, 715, 3900, 800, 0),
		(drawing, 3441, 716, 3900, 800, 0),
		(drawing, 3442, 716, 3900, 800, 0),
		(drawing, 3443, 716, 3900, 800, 0),
		(drawing, 3444, 716, 3900, 800, 0),
		(drawing, 3445, 716, 3900, 800, 0),
		(drawing, 3446, 716, 3900, 800, 0),
		(drawing, 3447, 717, 3900, 800, 0),
		(drawing, 3448, 717, 3900, 800, 0),
		(drawing, 3449, 717, 3900, 800, 0),
		(drawing, 3450, 717, 3900, 800, 0),
		(drawing, 3451, 717, 3900, 800, 0),
		(drawing, 3452, 718, 3900, 800, 0),
		(drawing, 3453, 718, 3900, 800, 0),
		(drawing, 3454, 718, 3900, 800, 0),
		(drawing, 3455, 718, 3900, 800, 0),
		(drawing, 3456, 718, 3900, 800, 0),
		(drawing, 3457, 719, 3900, 800, 0),
		(drawing, 3458, 719, 3900, 800, 0),
		(drawing, 3459, 719, 3900, 800, 0),
		(drawing, 3460, 719, 3900, 800, 0),
		(drawing, 3461, 719, 3900, 800, 0),
		(drawing, 3462, 719, 3900, 800, 0),
		(drawing, 3463, 720, 3900, 800, 0),
		(drawing, 3464, 720, 3900, 800, 0),
		(drawing, 3465, 720, 3900, 800, 0),
		(drawing, 3466, 720, 3900, 800, 0),
		(drawing, 3467, 720, 3900, 800, 0),
		(drawing, 3468, 721, 3900, 800, 0),
		(drawing, 3469, 721, 3900, 800, 0),
		(drawing, 3470, 721, 3900, 800, 0),
		(drawing, 3471, 721, 3900, 800, 0),
		(drawing, 3472, 721, 3900, 800, 0),
		(drawing, 3473, 721, 3900, 800, 0),
		(drawing, 3474, 722, 3900, 800, 0),
		(drawing, 3475, 722, 3900, 800, 0),
		(drawing, 3476, 722, 3900, 800, 0),
		(drawing, 3477, 722, 3900, 800, 0),
		(drawing, 3478, 722, 3900, 800, 0),
		(drawing, 3479, 723, 3900, 800, 0),
		(drawing, 3480, 723, 3900, 800, 0),
		(drawing, 3481, 723, 3900, 800, 0),
		(drawing, 3482, 723, 3900, 800, 0),
		(drawing, 3483, 723, 3900, 800, 0),
		(drawing, 3484, 723, 3900, 800, 0),
		(drawing, 3485, 724, 3900, 800, 0),
		(drawing, 3486, 724, 3900, 800, 0),
		(drawing, 3487, 724, 3900, 800, 0),
		(drawing, 3488, 724, 3900, 800, 0),
		(drawing, 3489, 724, 3900, 800, 0),
		(drawing, 3490, 725, 3900, 800, 0),
		(drawing, 3491, 725, 3900, 800, 0),
		(drawing, 3492, 725, 3900, 800, 0),
		(drawing, 3493, 725, 3900, 800, 0),
		(drawing, 3494, 725, 3900, 800, 0),
		(drawing, 3495, 725, 3900, 800, 0),
		(drawing, 3496, 726, 3900, 800, 0),
		(drawing, 3497, 726, 3900, 800, 0),
		(drawing, 3498, 726, 3900, 800, 0),
		(drawing, 3499, 726, 3900, 800, 0),
		(drawing, 3500, 726, 3900, 800, 0),
		(drawing, 3501, 727, 3900, 800, 0),
		(drawing, 3502, 727, 3900, 800, 0),
		(drawing, 3503, 727, 3900, 800, 0),
		(drawing, 3504, 727, 3900, 800, 0),
		(drawing, 3505, 727, 3900, 800, 0),
		(drawing, 3506, 728, 3900, 800, 0),
		(drawing, 3507, 728, 3900, 800, 0),
		(drawing, 3508, 728, 3900, 800, 0),
		(drawing, 3509, 728, 3900, 800, 0),
		(drawing, 3510, 728, 3900, 800, 0),
		(drawing, 3511, 728, 3900, 800, 0),
		(drawing, 3512, 729, 3900, 800, 0),
		(drawing, 3513, 729, 3900, 800, 0),
		(drawing, 3514, 729, 3900, 800, 0),
		(drawing, 3515, 729, 3900, 800, 0),
		(drawing, 3516, 729, 3900, 800, 0),
		(drawing, 3517, 730, 3900, 800, 0),
		(drawing, 3518, 730, 3900, 800, 0),
		(drawing, 3519, 730, 3900, 800, 0),
		(drawing, 3520, 730, 3900, 800, 0),
		(drawing, 3521, 730, 3900, 800, 0),
		(drawing, 3522, 730, 3900, 800, 0),
		(drawing, 3523, 731, 3900, 800, 0),
		(drawing, 3524, 731, 3900, 800, 0),
		(drawing, 3525, 731, 3900, 800, 0),
		(drawing, 3526, 731, 3900, 800, 0),
		(drawing, 3527, 731, 3900, 800, 0),
		(drawing, 3528, 732, 3900, 800, 0),
		(drawing, 3529, 732, 3900, 800, 0),
		(drawing, 3530, 732, 3900, 800, 0),
		(drawing, 3531, 732, 3900, 800, 0),
		(drawing, 3532, 732, 3900, 800, 0),
		(drawing, 3533, 732, 3900, 800, 0),
		(drawing, 3534, 733, 3900, 800, 0),
		(drawing, 3535, 733, 3900, 800, 0),
		(drawing, 3536, 733, 3900, 800, 0),
		(drawing, 3537, 733, 3900, 800, 0),
		(drawing, 3538, 733, 3900, 800, 0),
		(drawing, 3539, 734, 3900, 800, 0),
		(drawing, 3540, 734, 3900, 800, 0),
		(drawing, 3541, 734, 3900, 800, 0),
		(drawing, 3542, 734, 3900, 800, 0),
		(drawing, 3543, 734, 3900, 800, 0),
		(drawing, 3544, 735, 3900, 800, 0),
		(drawing, 3545, 735, 3900, 800, 0),
		(drawing, 3546, 735, 3900, 800, 0),
		(drawing, 3547, 735, 3900, 800, 0),
		(drawing, 3548, 735, 3900, 800, 0),
		(drawing, 3549, 735, 3900, 800, 0),
		(drawing, 3550, 736, 3900, 800, 0),
		(drawing, 3551, 736, 3900, 800, 0),
		(drawing, 3552, 736, 3900, 800, 0),
		(drawing, 3553, 736, 3900, 800, 0),
		(drawing, 3554, 736, 3900, 800, 0),
		(drawing, 3555, 737, 3900, 800, 0),
		(drawing, 3556, 737, 3900, 800, 0),
		(drawing, 3557, 737, 3900, 800, 0),
		(drawing, 3558, 737, 3900, 800, 0),
		(drawing, 3559, 737, 3900, 800, 0),
		(drawing, 3560, 737, 3900, 800, 0),
		(drawing, 3561, 738, 3900, 800, 0),
		(drawing, 3562, 738, 3900, 800, 0),
		(drawing, 3563, 738, 3900, 800, 0),
		(drawing, 3564, 738, 3900, 800, 0),
		(drawing, 3565, 738, 3900, 800, 0),
		(drawing, 3566, 739, 3900, 800, 0),
		(drawing, 3567, 739, 3900, 800, 0),
		(drawing, 3568, 739, 3900, 800, 0),
		(drawing, 3569, 739, 3900, 800, 0),
		(drawing, 3570, 739, 3900, 800, 0),
		(drawing, 3571, 739, 3900, 800, 0),
		(drawing, 3572, 740, 3900, 800, 0),
		(drawing, 3573, 740, 3900, 800, 0),
		(drawing, 3574, 740, 3900, 800, 0),
		(drawing, 3575, 740, 3900, 800, 0),
		(drawing, 3576, 740, 3900, 800, 0),
		(drawing, 3577, 741, 3900, 800, 0),
		(drawing, 3578, 741, 3900, 800, 0),
		(drawing, 3579, 741, 3900, 800, 0),
		(drawing, 3580, 741, 3900, 800, 0),
		(drawing, 3581, 741, 3900, 800, 0),
		(drawing, 3582, 742, 3900, 800, 0),
		(drawing, 3583, 742, 3900, 800, 0),
		(drawing, 3584, 742, 3900, 800, 0),
		(drawing, 3585, 742, 3900, 800, 0),
		(drawing, 3586, 742, 3900, 800, 0),
		(drawing, 3587, 742, 3900, 800, 0),
		(drawing, 3588, 743, 3900, 800, 0),
		(drawing, 3589, 743, 3900, 800, 0),
		(drawing, 3590, 743, 3900, 800, 0),
		(drawing, 3591, 743, 3900, 800, 0),
		(drawing, 3592, 743, 3900, 800, 0),
		(drawing, 3593, 744, 3900, 800, 0),
		(drawing, 3594, 744, 3900, 800, 0),
		(drawing, 3595, 744, 3900, 800, 0),
		(drawing, 3596, 744, 3900, 800, 0),
		(drawing, 3597, 744, 3900, 800, 0),
		(drawing, 3598, 744, 3900, 800, 0),
		(drawing, 3599, 745, 3900, 800, 0),
		(drawing, 3600, 745, 3900, 800, 0),
		(drawing, 3601, 745, 3900, 800, 0),
		(drawing, 3602, 745, 3900, 800, 0),
		(drawing, 3603, 745, 3900, 800, 0),
		(drawing, 3604, 746, 3900, 800, 0),
		(drawing, 3605, 746, 3900, 800, 0),
		(drawing, 3606, 746, 3900, 800, 0),
		(drawing, 3607, 746, 3900, 800, 0),
		(drawing, 3608, 746, 3900, 800, 0),
		(drawing, 3609, 746, 3900, 800, 0),
		(drawing, 3610, 747, 3900, 800, 0),
		(drawing, 3611, 747, 3900, 800, 0),
		(drawing, 3612, 747, 3900, 800, 0),
		(drawing, 3613, 747, 3900, 800, 0),
		(drawing, 3614, 747, 3900, 800, 0),
		(drawing, 3615, 748, 3900, 800, 0),
		(drawing, 3616, 748, 3900, 800, 0),
		(drawing, 3617, 748, 3900, 800, 0),
		(drawing, 3618, 748, 3900, 800, 0),
		(drawing, 3619, 748, 3900, 800, 0),
		(drawing, 3620, 748, 3900, 800, 0),
		(drawing, 3621, 749, 3900, 800, 0),
		(drawing, 3622, 749, 3900, 800, 0),
		(drawing, 3623, 749, 3900, 800, 0),
		(drawing, 3624, 749, 3900, 800, 0),
		(drawing, 3625, 749, 3900, 800, 0),
		(drawing, 3626, 750, 3900, 800, 0),
		(drawing, 3627, 750, 3900, 800, 0),
		(drawing, 3628, 750, 3900, 800, 0),
		(drawing, 3629, 750, 3900, 800, 0),
		(drawing, 3630, 750, 3900, 800, 0),
		(drawing, 3631, 751, 3900, 800, 0),
		(drawing, 3632, 751, 3900, 800, 0),
		(drawing, 3633, 751, 3900, 800, 0),
		(drawing, 3634, 751, 3900, 800, 0),
		(drawing, 3635, 751, 3900, 800, 0),
		(drawing, 3636, 751, 3900, 800, 0),
		(drawing, 3637, 752, 3900, 800, 0),
		(drawing, 3638, 752, 3900, 800, 0),
		(drawing, 3639, 752, 3900, 800, 0),
		(drawing, 3640, 752, 3900, 800, 0),
		(drawing, 3641, 752, 3900, 800, 0),
		(drawing, 3642, 753, 3900, 800, 0),
		(drawing, 3643, 753, 3900, 800, 0),
		(drawing, 3644, 753, 3900, 800, 0),
		(drawing, 3645, 753, 3900, 800, 0),
		(drawing, 3646, 753, 3900, 800, 0),
		(drawing, 3647, 753, 3900, 800, 0),
		(drawing, 3648, 754, 3900, 800, 0),
		(drawing, 3649, 754, 3900, 800, 0),
		(drawing, 3650, 754, 3900, 800, 0),
		(drawing, 3651, 754, 3900, 800, 0),
		(drawing, 3652, 754, 3900, 800, 0),
		(drawing, 3653, 755, 3900, 800, 0),
		(drawing, 3654, 755, 3900, 800, 0),
		(drawing, 3655, 755, 3900, 800, 0),
		(drawing, 3656, 755, 3900, 800, 0),
		(drawing, 3657, 755, 3900, 800, 0),
		(drawing, 3658, 755, 3900, 800, 0),
		(drawing, 3659, 756, 3900, 800, 0),
		(drawing, 3660, 756, 3900, 800, 0),
		(drawing, 3661, 756, 3900, 800, 0),
		(drawing, 3662, 756, 3900, 800, 0),
		(drawing, 3663, 756, 3900, 800, 0),
		(drawing, 3664, 757, 3900, 800, 0),
		(drawing, 3665, 757, 3900, 800, 0),
		(drawing, 3666, 757, 3900, 800, 0),
		(drawing, 3667, 757, 3900, 800, 0),
		(drawing, 3668, 757, 3900, 800, 0),
		(drawing, 3669, 758, 3900, 800, 0),
		(drawing, 3670, 758, 3900, 800, 0),
		(drawing, 3671, 758, 3900, 800, 0),
		(drawing, 3672, 758, 3900, 800, 0),
		(drawing, 3673, 758, 3900, 800, 0),
		(drawing, 3674, 758, 3900, 800, 0),
		(drawing, 3675, 759, 3900, 800, 0),
		(drawing, 3676, 759, 3900, 800, 0),
		(drawing, 3677, 759, 3900, 800, 0),
		(drawing, 3678, 759, 3900, 800, 0),
		(drawing, 3679, 759, 3900, 800, 0),
		(drawing, 3680, 760, 3900, 800, 0),
		(drawing, 3681, 760, 3900, 800, 0),
		(drawing, 3682, 760, 3900, 800, 0),
		(drawing, 3683, 760, 3900, 800, 0),
		(drawing, 3684, 760, 3900, 800, 0),
		(drawing, 3685, 760, 3900, 800, 0),
		(drawing, 3686, 761, 3900, 800, 0),
		(drawing, 3687, 761, 3900, 800, 0),
		(drawing, 3688, 761, 3900, 800, 0),
		(drawing, 3689, 761, 3900, 800, 0),
		(drawing, 3690, 761, 3900, 800, 0),
		(drawing, 3691, 762, 3900, 800, 0),
		(drawing, 3692, 762, 3900, 800, 0),
		(drawing, 3693, 762, 3900, 800, 0),
		(drawing, 3694, 762, 3900, 800, 0),
		(drawing, 3695, 762, 3900, 800, 0),
		(drawing, 3696, 762, 3900, 800, 0),
		(drawing, 3697, 763, 3900, 800, 0),
		(drawing, 3698, 763, 3900, 800, 0),
		(drawing, 3699, 763, 3900, 800, 0),
		(drawing, 3700, 763, 3900, 800, 0),
		(drawing, 3701, 763, 3900, 800, 0),
		(drawing, 3702, 764, 3900, 800, 0),
		(drawing, 3703, 764, 3900, 800, 0),
		(drawing, 3704, 764, 3900, 800, 0),
		(drawing, 3705, 764, 3900, 800, 0),
		(drawing, 3706, 764, 3900, 800, 0),
		(drawing, 3707, 764, 3900, 800, 0),
		(drawing, 3708, 765, 3900, 800, 0),
		(drawing, 3709, 765, 3900, 800, 0),
		(drawing, 3710, 765, 3900, 800, 0),
		(drawing, 3711, 765, 3900, 800, 0),
		(drawing, 3712, 765, 3900, 800, 0),
		(drawing, 3713, 766, 3900, 800, 0),
		(drawing, 3714, 766, 3900, 800, 0),
		(drawing, 3715, 766, 3900, 800, 0),
		(drawing, 3716, 766, 3900, 800, 0),
		(drawing, 3717, 766, 3900, 800, 0),
		(drawing, 3718, 767, 3900, 800, 0),
		(drawing, 3719, 767, 3900, 800, 0),
		(drawing, 3720, 767, 3900, 800, 0),
		(drawing, 3721, 767, 3900, 800, 0),
		(drawing, 3722, 767, 3900, 800, 0),
		(drawing, 3723, 767, 3900, 800, 0),
		(drawing, 3724, 768, 3900, 800, 0),
		(drawing, 3725, 768, 3900, 800, 0),
		(drawing, 3726, 768, 3900, 800, 0),
		(drawing, 3727, 768, 3900, 800, 0),
		(drawing, 3728, 768, 3900, 800, 0),
		(drawing, 3729, 769, 3900, 800, 0),
		(drawing, 3730, 769, 3900, 800, 0),
		(drawing, 3731, 769, 3900, 800, 0),
		(drawing, 3732, 769, 3900, 800, 0),
		(drawing, 3733, 769, 3900, 800, 0),
		(drawing, 3734, 769, 3900, 800, 0),
		(drawing, 3735, 770, 3900, 800, 0),
		(drawing, 3736, 770, 3900, 800, 0),
		(drawing, 3737, 770, 3900, 800, 0),
		(drawing, 3738, 770, 3900, 800, 0),
		(drawing, 3739, 770, 3900, 800, 0),
		(drawing, 3740, 771, 3900, 800, 0),
		(drawing, 3741, 771, 3900, 800, 0),
		(drawing, 3742, 771, 3900, 800, 0),
		(drawing, 3743, 771, 3900, 800, 0),
		(drawing, 3744, 771, 3900, 800, 0),
		(drawing, 3745, 771, 3900, 800, 0),
		(drawing, 3746, 772, 3900, 800, 0),
		(drawing, 3747, 772, 3900, 800, 0),
		(drawing, 3748, 772, 3900, 800, 0),
		(drawing, 3749, 772, 3900, 800, 0),
		(drawing, 3750, 772, 3900, 800, 0),
		(drawing, 3751, 773, 3900, 800, 0),
		(drawing, 3752, 773, 3900, 800, 0),
		(drawing, 3753, 773, 3900, 800, 0),
		(drawing, 3754, 773, 3900, 800, 0),
		(drawing, 3755, 773, 3900, 800, 0),
		(drawing, 3756, 774, 3900, 800, 0),
		(drawing, 3757, 774, 3900, 800, 0),
		(drawing, 3758, 774, 3900, 800, 0),
		(drawing, 3759, 774, 3900, 800, 0),
		(drawing, 3760, 774, 3900, 800, 0),
		(drawing, 3761, 774, 3900, 800, 0),
		(drawing, 3762, 775, 3900, 800, 0),
		(drawing, 3763, 775, 3900, 800, 0),
		(drawing, 3764, 775, 3900, 800, 0),
		(drawing, 3765, 775, 3900, 800, 0),
		(drawing, 3766, 775, 3900, 800, 0),
		(drawing, 3767, 776, 3900, 800, 0),
		(drawing, 3768, 776, 3900, 800, 0),
		(drawing, 3769, 776, 3900, 800, 0),
		(drawing, 3770, 776, 3900, 800, 0),
		(drawing, 3771, 776, 3900, 800, 0),
		(drawing, 3772, 776, 3900, 800, 0),
		(drawing, 3773, 777, 3900, 800, 0),
		(drawing, 3774, 777, 3900, 800, 0),
		(drawing, 3775, 777, 3900, 800, 0),
		(drawing, 3776, 777, 3900, 800, 0),
		(drawing, 3777, 777, 3900, 800, 0),
		(drawing, 3778, 778, 3900, 800, 0),
		(drawing, 3779, 778, 3900, 800, 0),
		(drawing, 3780, 778, 3900, 800, 0),
		(drawing, 3781, 778, 3900, 800, 0),
		(drawing, 3782, 778, 3900, 800, 0),
		(drawing, 3783, 778, 3900, 800, 0),
		(drawing, 3784, 779, 3900, 800, 0),
		(drawing, 3785, 779, 3900, 800, 0),
		(drawing, 3786, 779, 3900, 800, 0),
		(drawing, 3787, 779, 3900, 800, 0),
		(drawing, 3788, 779, 3900, 800, 0),
		(drawing, 3789, 780, 3900, 800, 0),
		(drawing, 3790, 780, 3900, 800, 0),
		(drawing, 3791, 780, 3900, 800, 0),
		(drawing, 3792, 780, 3900, 800, 0),
		(drawing, 3793, 780, 3900, 800, 0),
		(drawing, 3794, 781, 3900, 800, 0),
		(drawing, 3795, 781, 3900, 800, 0),
		(drawing, 3796, 781, 3900, 800, 0),
		(drawing, 3797, 781, 3900, 800, 0),
		(drawing, 3798, 781, 3900, 800, 0),
		(drawing, 3799, 781, 3900, 800, 0),
		(drawing, 3800, 782, 3900, 800, 0),
		(drawing, 3801, 782, 3900, 800, 0),
		(drawing, 3802, 782, 3900, 800, 0),
		(drawing, 3803, 782, 3900, 800, 0),
		(drawing, 3804, 782, 3900, 800, 0),
		(drawing, 3805, 783, 3900, 800, 0),
		(drawing, 3806, 783, 3900, 800, 0),
		(drawing, 3807, 783, 3900, 800, 0),
		(drawing, 3808, 783, 3900, 800, 0),
		(drawing, 3809, 783, 3900, 800, 0),
		(drawing, 3810, 783, 3900, 800, 0),
		(drawing, 3811, 784, 3900, 800, 0),
		(drawing, 3812, 784, 3900, 800, 0),
		(drawing, 3813, 784, 3900, 800, 0),
		(drawing, 3814, 784, 3900, 800, 0),
		(drawing, 3815, 784, 3900, 800, 0),
		(drawing, 3816, 785, 3900, 800, 0),
		(drawing, 3817, 785, 3900, 800, 0),
		(drawing, 3818, 785, 3900, 800, 0),
		(drawing, 3819, 785, 3900, 800, 0),
		(drawing, 3820, 785, 3900, 800, 0),
		(drawing, 3821, 785, 3900, 800, 0),
		(drawing, 3822, 786, 3900, 800, 0),
		(drawing, 3823, 786, 3900, 800, 0),
		(drawing, 3824, 786, 3900, 800, 0),
		(drawing, 3825, 786, 3900, 800, 0),
		(drawing, 3826, 786, 3900, 800, 0),
		(drawing, 3827, 787, 3900, 800, 0),
		(drawing, 3828, 787, 3900, 800, 0),
		(drawing, 3829, 787, 3900, 800, 0),
		(drawing, 3830, 787, 3900, 800, 0),
		(drawing, 3831, 787, 3900, 800, 0),
		(drawing, 3832, 787, 3900, 800, 0),
		(drawing, 3833, 788, 3900, 800, 0),
		(drawing, 3834, 788, 3900, 800, 0),
		(drawing, 3835, 788, 3900, 800, 0),
		(drawing, 3836, 788, 3900, 800, 0),
		(drawing, 3837, 788, 3900, 800, 0),
		(drawing, 3838, 789, 3900, 800, 0),
		(drawing, 3839, 789, 3900, 800, 0),
		(drawing, 3840, 789, 3900, 800, 0),
		(drawing, 3841, 789, 3900, 800, 0),
		(drawing, 3842, 789, 3900, 800, 0),
		(drawing, 3843, 790, 3900, 800, 0),
		(drawing, 3844, 790, 3900, 800, 0),
		(drawing, 3845, 790, 3900, 800, 0),
		(drawing, 3846, 790, 3900, 800, 0),
		(drawing, 3847, 790, 3900, 800, 0),
		(drawing, 3848, 790, 3900, 800, 0),
		(drawing, 3849, 791, 3900, 800, 0),
		(drawing, 3850, 791, 3900, 800, 0),
		(drawing, 3851, 791, 3900, 800, 0),
		(drawing, 3852, 791, 3900, 800, 0),
		(drawing, 3853, 791, 3900, 800, 0),
		(drawing, 3854, 792, 3900, 800, 0),
		(drawing, 3855, 792, 3900, 800, 0),
		(drawing, 3856, 792, 3900, 800, 0),
		(drawing, 3857, 792, 3900, 800, 0),
		(drawing, 3858, 792, 3900, 800, 0),
		(drawing, 3859, 792, 3900, 800, 0),
		(drawing, 3860, 793, 3900, 800, 0),
		(drawing, 3861, 793, 3900, 800, 0),
		(drawing, 3862, 793, 3900, 800, 0),
		(drawing, 3863, 793, 3900, 800, 0),
		(drawing, 3864, 793, 3900, 800, 0),
		(drawing, 3865, 794, 3900, 800, 0),
		(drawing, 3866, 794, 3900, 800, 0),
		(drawing, 3867, 794, 3900, 800, 0),
		(drawing, 3868, 794, 3900, 800, 0),
		(drawing, 3869, 794, 3900, 800, 0),
		(drawing, 3870, 794, 3900, 800, 0),
		(drawing, 3871, 795, 3900, 800, 0),
		(drawing, 3872, 795, 3900, 800, 0),
		(drawing, 3873, 795, 3900, 800, 0),
		(drawing, 3874, 795, 3900, 800, 0),
		(drawing, 3875, 795, 3900, 800, 0),
		(drawing, 3876, 796, 3900, 800, 0),
		(drawing, 3877, 796, 3900, 800, 0),
		(drawing, 3878, 796, 3900, 800, 0),
		(drawing, 3879, 796, 3900, 800, 0),
		(drawing, 3880, 796, 3900, 800, 0),
		(drawing, 3881, 797, 3900, 800, 0),
		(drawing, 3882, 797, 3900, 800, 0),
		(drawing, 3883, 797, 3900, 800, 0),
		(drawing, 3884, 797, 3900, 800, 0),
		(drawing, 3885, 797, 3900, 800, 0),
		(drawing, 3886, 797, 3900, 800, 0),
		(drawing, 3887, 798, 3900, 800, 0),
		(drawing, 3888, 798, 3900, 800, 0),
		(drawing, 3889, 798, 3900, 800, 0),
		(drawing, 3890, 798, 3900, 800, 0),
		(drawing, 3891, 798, 3900, 800, 0),
		(drawing, 3892, 799, 3900, 800, 0),
		(drawing, 3893, 799, 3900, 800, 0),
		(drawing, 3894, 799, 3900, 800, 0),
		(drawing, 3895, 799, 3900, 800, 0),
		(drawing, 3896, 799, 3900, 800, 0),
		(drawing, 3897, 799, 3900, 800, 0),
		(drawing, 3898, 800, 3900, 800, 0),
		(drawing, 3899, 800, 3900, 800, 0),
		(done, 3900, 800, 3900, 800, 0)
	);
END PACKAGE ex1_data_pak;
