-- advanced test 3
-- draw line from (0,0) to (4095,0)
-- NOTE * xincr is a 12bits logic vector
--------* the maximum value of it is b1111,1111,1111 which is 4095 in decimal
--------* this test is for the case of maximum possible value of xincr

PACKAGE ex1_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 0, 0, 0),
		(start, 0, 0, 4095, 0, 0),
		(drawing, 0, 0, 4095, 0, 0),
		(drawing, 1, 0, 4095, 0, 0),
		(drawing, 2, 0, 4095, 0, 0),
		(drawing, 3, 0, 4095, 0, 0),
		(drawing, 4, 0, 4095, 0, 0),
		(drawing, 5, 0, 4095, 0, 0),
		(drawing, 6, 0, 4095, 0, 0),
		(drawing, 7, 0, 4095, 0, 0),
		(drawing, 8, 0, 4095, 0, 0),
		(drawing, 9, 0, 4095, 0, 0),
		(drawing, 10, 0, 4095, 0, 0),
		(drawing, 11, 0, 4095, 0, 0),
		(drawing, 12, 0, 4095, 0, 0),
		(drawing, 13, 0, 4095, 0, 0),
		(drawing, 14, 0, 4095, 0, 0),
		(drawing, 15, 0, 4095, 0, 0),
		(drawing, 16, 0, 4095, 0, 0),
		(drawing, 17, 0, 4095, 0, 0),
		(drawing, 18, 0, 4095, 0, 0),
		(drawing, 19, 0, 4095, 0, 0),
		(drawing, 20, 0, 4095, 0, 0),
		(drawing, 21, 0, 4095, 0, 0),
		(drawing, 22, 0, 4095, 0, 0),
		(drawing, 23, 0, 4095, 0, 0),
		(drawing, 24, 0, 4095, 0, 0),
		(drawing, 25, 0, 4095, 0, 0),
		(drawing, 26, 0, 4095, 0, 0),
		(drawing, 27, 0, 4095, 0, 0),
		(drawing, 28, 0, 4095, 0, 0),
		(drawing, 29, 0, 4095, 0, 0),
		(drawing, 30, 0, 4095, 0, 0),
		(drawing, 31, 0, 4095, 0, 0),
		(drawing, 32, 0, 4095, 0, 0),
		(drawing, 33, 0, 4095, 0, 0),
		(drawing, 34, 0, 4095, 0, 0),
		(drawing, 35, 0, 4095, 0, 0),
		(drawing, 36, 0, 4095, 0, 0),
		(drawing, 37, 0, 4095, 0, 0),
		(drawing, 38, 0, 4095, 0, 0),
		(drawing, 39, 0, 4095, 0, 0),
		(drawing, 40, 0, 4095, 0, 0),
		(drawing, 41, 0, 4095, 0, 0),
		(drawing, 42, 0, 4095, 0, 0),
		(drawing, 43, 0, 4095, 0, 0),
		(drawing, 44, 0, 4095, 0, 0),
		(drawing, 45, 0, 4095, 0, 0),
		(drawing, 46, 0, 4095, 0, 0),
		(drawing, 47, 0, 4095, 0, 0),
		(drawing, 48, 0, 4095, 0, 0),
		(drawing, 49, 0, 4095, 0, 0),
		(drawing, 50, 0, 4095, 0, 0),
		(drawing, 51, 0, 4095, 0, 0),
		(drawing, 52, 0, 4095, 0, 0),
		(drawing, 53, 0, 4095, 0, 0),
		(drawing, 54, 0, 4095, 0, 0),
		(drawing, 55, 0, 4095, 0, 0),
		(drawing, 56, 0, 4095, 0, 0),
		(drawing, 57, 0, 4095, 0, 0),
		(drawing, 58, 0, 4095, 0, 0),
		(drawing, 59, 0, 4095, 0, 0),
		(drawing, 60, 0, 4095, 0, 0),
		(drawing, 61, 0, 4095, 0, 0),
		(drawing, 62, 0, 4095, 0, 0),
		(drawing, 63, 0, 4095, 0, 0),
		(drawing, 64, 0, 4095, 0, 0),
		(drawing, 65, 0, 4095, 0, 0),
		(drawing, 66, 0, 4095, 0, 0),
		(drawing, 67, 0, 4095, 0, 0),
		(drawing, 68, 0, 4095, 0, 0),
		(drawing, 69, 0, 4095, 0, 0),
		(drawing, 70, 0, 4095, 0, 0),
		(drawing, 71, 0, 4095, 0, 0),
		(drawing, 72, 0, 4095, 0, 0),
		(drawing, 73, 0, 4095, 0, 0),
		(drawing, 74, 0, 4095, 0, 0),
		(drawing, 75, 0, 4095, 0, 0),
		(drawing, 76, 0, 4095, 0, 0),
		(drawing, 77, 0, 4095, 0, 0),
		(drawing, 78, 0, 4095, 0, 0),
		(drawing, 79, 0, 4095, 0, 0),
		(drawing, 80, 0, 4095, 0, 0),
		(drawing, 81, 0, 4095, 0, 0),
		(drawing, 82, 0, 4095, 0, 0),
		(drawing, 83, 0, 4095, 0, 0),
		(drawing, 84, 0, 4095, 0, 0),
		(drawing, 85, 0, 4095, 0, 0),
		(drawing, 86, 0, 4095, 0, 0),
		(drawing, 87, 0, 4095, 0, 0),
		(drawing, 88, 0, 4095, 0, 0),
		(drawing, 89, 0, 4095, 0, 0),
		(drawing, 90, 0, 4095, 0, 0),
		(drawing, 91, 0, 4095, 0, 0),
		(drawing, 92, 0, 4095, 0, 0),
		(drawing, 93, 0, 4095, 0, 0),
		(drawing, 94, 0, 4095, 0, 0),
		(drawing, 95, 0, 4095, 0, 0),
		(drawing, 96, 0, 4095, 0, 0),
		(drawing, 97, 0, 4095, 0, 0),
		(drawing, 98, 0, 4095, 0, 0),
		(drawing, 99, 0, 4095, 0, 0),
		(drawing, 100, 0, 4095, 0, 0),
		(drawing, 101, 0, 4095, 0, 0),
		(drawing, 102, 0, 4095, 0, 0),
		(drawing, 103, 0, 4095, 0, 0),
		(drawing, 104, 0, 4095, 0, 0),
		(drawing, 105, 0, 4095, 0, 0),
		(drawing, 106, 0, 4095, 0, 0),
		(drawing, 107, 0, 4095, 0, 0),
		(drawing, 108, 0, 4095, 0, 0),
		(drawing, 109, 0, 4095, 0, 0),
		(drawing, 110, 0, 4095, 0, 0),
		(drawing, 111, 0, 4095, 0, 0),
		(drawing, 112, 0, 4095, 0, 0),
		(drawing, 113, 0, 4095, 0, 0),
		(drawing, 114, 0, 4095, 0, 0),
		(drawing, 115, 0, 4095, 0, 0),
		(drawing, 116, 0, 4095, 0, 0),
		(drawing, 117, 0, 4095, 0, 0),
		(drawing, 118, 0, 4095, 0, 0),
		(drawing, 119, 0, 4095, 0, 0),
		(drawing, 120, 0, 4095, 0, 0),
		(drawing, 121, 0, 4095, 0, 0),
		(drawing, 122, 0, 4095, 0, 0),
		(drawing, 123, 0, 4095, 0, 0),
		(drawing, 124, 0, 4095, 0, 0),
		(drawing, 125, 0, 4095, 0, 0),
		(drawing, 126, 0, 4095, 0, 0),
		(drawing, 127, 0, 4095, 0, 0),
		(drawing, 128, 0, 4095, 0, 0),
		(drawing, 129, 0, 4095, 0, 0),
		(drawing, 130, 0, 4095, 0, 0),
		(drawing, 131, 0, 4095, 0, 0),
		(drawing, 132, 0, 4095, 0, 0),
		(drawing, 133, 0, 4095, 0, 0),
		(drawing, 134, 0, 4095, 0, 0),
		(drawing, 135, 0, 4095, 0, 0),
		(drawing, 136, 0, 4095, 0, 0),
		(drawing, 137, 0, 4095, 0, 0),
		(drawing, 138, 0, 4095, 0, 0),
		(drawing, 139, 0, 4095, 0, 0),
		(drawing, 140, 0, 4095, 0, 0),
		(drawing, 141, 0, 4095, 0, 0),
		(drawing, 142, 0, 4095, 0, 0),
		(drawing, 143, 0, 4095, 0, 0),
		(drawing, 144, 0, 4095, 0, 0),
		(drawing, 145, 0, 4095, 0, 0),
		(drawing, 146, 0, 4095, 0, 0),
		(drawing, 147, 0, 4095, 0, 0),
		(drawing, 148, 0, 4095, 0, 0),
		(drawing, 149, 0, 4095, 0, 0),
		(drawing, 150, 0, 4095, 0, 0),
		(drawing, 151, 0, 4095, 0, 0),
		(drawing, 152, 0, 4095, 0, 0),
		(drawing, 153, 0, 4095, 0, 0),
		(drawing, 154, 0, 4095, 0, 0),
		(drawing, 155, 0, 4095, 0, 0),
		(drawing, 156, 0, 4095, 0, 0),
		(drawing, 157, 0, 4095, 0, 0),
		(drawing, 158, 0, 4095, 0, 0),
		(drawing, 159, 0, 4095, 0, 0),
		(drawing, 160, 0, 4095, 0, 0),
		(drawing, 161, 0, 4095, 0, 0),
		(drawing, 162, 0, 4095, 0, 0),
		(drawing, 163, 0, 4095, 0, 0),
		(drawing, 164, 0, 4095, 0, 0),
		(drawing, 165, 0, 4095, 0, 0),
		(drawing, 166, 0, 4095, 0, 0),
		(drawing, 167, 0, 4095, 0, 0),
		(drawing, 168, 0, 4095, 0, 0),
		(drawing, 169, 0, 4095, 0, 0),
		(drawing, 170, 0, 4095, 0, 0),
		(drawing, 171, 0, 4095, 0, 0),
		(drawing, 172, 0, 4095, 0, 0),
		(drawing, 173, 0, 4095, 0, 0),
		(drawing, 174, 0, 4095, 0, 0),
		(drawing, 175, 0, 4095, 0, 0),
		(drawing, 176, 0, 4095, 0, 0),
		(drawing, 177, 0, 4095, 0, 0),
		(drawing, 178, 0, 4095, 0, 0),
		(drawing, 179, 0, 4095, 0, 0),
		(drawing, 180, 0, 4095, 0, 0),
		(drawing, 181, 0, 4095, 0, 0),
		(drawing, 182, 0, 4095, 0, 0),
		(drawing, 183, 0, 4095, 0, 0),
		(drawing, 184, 0, 4095, 0, 0),
		(drawing, 185, 0, 4095, 0, 0),
		(drawing, 186, 0, 4095, 0, 0),
		(drawing, 187, 0, 4095, 0, 0),
		(drawing, 188, 0, 4095, 0, 0),
		(drawing, 189, 0, 4095, 0, 0),
		(drawing, 190, 0, 4095, 0, 0),
		(drawing, 191, 0, 4095, 0, 0),
		(drawing, 192, 0, 4095, 0, 0),
		(drawing, 193, 0, 4095, 0, 0),
		(drawing, 194, 0, 4095, 0, 0),
		(drawing, 195, 0, 4095, 0, 0),
		(drawing, 196, 0, 4095, 0, 0),
		(drawing, 197, 0, 4095, 0, 0),
		(drawing, 198, 0, 4095, 0, 0),
		(drawing, 199, 0, 4095, 0, 0),
		(drawing, 200, 0, 4095, 0, 0),
		(drawing, 201, 0, 4095, 0, 0),
		(drawing, 202, 0, 4095, 0, 0),
		(drawing, 203, 0, 4095, 0, 0),
		(drawing, 204, 0, 4095, 0, 0),
		(drawing, 205, 0, 4095, 0, 0),
		(drawing, 206, 0, 4095, 0, 0),
		(drawing, 207, 0, 4095, 0, 0),
		(drawing, 208, 0, 4095, 0, 0),
		(drawing, 209, 0, 4095, 0, 0),
		(drawing, 210, 0, 4095, 0, 0),
		(drawing, 211, 0, 4095, 0, 0),
		(drawing, 212, 0, 4095, 0, 0),
		(drawing, 213, 0, 4095, 0, 0),
		(drawing, 214, 0, 4095, 0, 0),
		(drawing, 215, 0, 4095, 0, 0),
		(drawing, 216, 0, 4095, 0, 0),
		(drawing, 217, 0, 4095, 0, 0),
		(drawing, 218, 0, 4095, 0, 0),
		(drawing, 219, 0, 4095, 0, 0),
		(drawing, 220, 0, 4095, 0, 0),
		(drawing, 221, 0, 4095, 0, 0),
		(drawing, 222, 0, 4095, 0, 0),
		(drawing, 223, 0, 4095, 0, 0),
		(drawing, 224, 0, 4095, 0, 0),
		(drawing, 225, 0, 4095, 0, 0),
		(drawing, 226, 0, 4095, 0, 0),
		(drawing, 227, 0, 4095, 0, 0),
		(drawing, 228, 0, 4095, 0, 0),
		(drawing, 229, 0, 4095, 0, 0),
		(drawing, 230, 0, 4095, 0, 0),
		(drawing, 231, 0, 4095, 0, 0),
		(drawing, 232, 0, 4095, 0, 0),
		(drawing, 233, 0, 4095, 0, 0),
		(drawing, 234, 0, 4095, 0, 0),
		(drawing, 235, 0, 4095, 0, 0),
		(drawing, 236, 0, 4095, 0, 0),
		(drawing, 237, 0, 4095, 0, 0),
		(drawing, 238, 0, 4095, 0, 0),
		(drawing, 239, 0, 4095, 0, 0),
		(drawing, 240, 0, 4095, 0, 0),
		(drawing, 241, 0, 4095, 0, 0),
		(drawing, 242, 0, 4095, 0, 0),
		(drawing, 243, 0, 4095, 0, 0),
		(drawing, 244, 0, 4095, 0, 0),
		(drawing, 245, 0, 4095, 0, 0),
		(drawing, 246, 0, 4095, 0, 0),
		(drawing, 247, 0, 4095, 0, 0),
		(drawing, 248, 0, 4095, 0, 0),
		(drawing, 249, 0, 4095, 0, 0),
		(drawing, 250, 0, 4095, 0, 0),
		(drawing, 251, 0, 4095, 0, 0),
		(drawing, 252, 0, 4095, 0, 0),
		(drawing, 253, 0, 4095, 0, 0),
		(drawing, 254, 0, 4095, 0, 0),
		(drawing, 255, 0, 4095, 0, 0),
		(drawing, 256, 0, 4095, 0, 0),
		(drawing, 257, 0, 4095, 0, 0),
		(drawing, 258, 0, 4095, 0, 0),
		(drawing, 259, 0, 4095, 0, 0),
		(drawing, 260, 0, 4095, 0, 0),
		(drawing, 261, 0, 4095, 0, 0),
		(drawing, 262, 0, 4095, 0, 0),
		(drawing, 263, 0, 4095, 0, 0),
		(drawing, 264, 0, 4095, 0, 0),
		(drawing, 265, 0, 4095, 0, 0),
		(drawing, 266, 0, 4095, 0, 0),
		(drawing, 267, 0, 4095, 0, 0),
		(drawing, 268, 0, 4095, 0, 0),
		(drawing, 269, 0, 4095, 0, 0),
		(drawing, 270, 0, 4095, 0, 0),
		(drawing, 271, 0, 4095, 0, 0),
		(drawing, 272, 0, 4095, 0, 0),
		(drawing, 273, 0, 4095, 0, 0),
		(drawing, 274, 0, 4095, 0, 0),
		(drawing, 275, 0, 4095, 0, 0),
		(drawing, 276, 0, 4095, 0, 0),
		(drawing, 277, 0, 4095, 0, 0),
		(drawing, 278, 0, 4095, 0, 0),
		(drawing, 279, 0, 4095, 0, 0),
		(drawing, 280, 0, 4095, 0, 0),
		(drawing, 281, 0, 4095, 0, 0),
		(drawing, 282, 0, 4095, 0, 0),
		(drawing, 283, 0, 4095, 0, 0),
		(drawing, 284, 0, 4095, 0, 0),
		(drawing, 285, 0, 4095, 0, 0),
		(drawing, 286, 0, 4095, 0, 0),
		(drawing, 287, 0, 4095, 0, 0),
		(drawing, 288, 0, 4095, 0, 0),
		(drawing, 289, 0, 4095, 0, 0),
		(drawing, 290, 0, 4095, 0, 0),
		(drawing, 291, 0, 4095, 0, 0),
		(drawing, 292, 0, 4095, 0, 0),
		(drawing, 293, 0, 4095, 0, 0),
		(drawing, 294, 0, 4095, 0, 0),
		(drawing, 295, 0, 4095, 0, 0),
		(drawing, 296, 0, 4095, 0, 0),
		(drawing, 297, 0, 4095, 0, 0),
		(drawing, 298, 0, 4095, 0, 0),
		(drawing, 299, 0, 4095, 0, 0),
		(drawing, 300, 0, 4095, 0, 0),
		(drawing, 301, 0, 4095, 0, 0),
		(drawing, 302, 0, 4095, 0, 0),
		(drawing, 303, 0, 4095, 0, 0),
		(drawing, 304, 0, 4095, 0, 0),
		(drawing, 305, 0, 4095, 0, 0),
		(drawing, 306, 0, 4095, 0, 0),
		(drawing, 307, 0, 4095, 0, 0),
		(drawing, 308, 0, 4095, 0, 0),
		(drawing, 309, 0, 4095, 0, 0),
		(drawing, 310, 0, 4095, 0, 0),
		(drawing, 311, 0, 4095, 0, 0),
		(drawing, 312, 0, 4095, 0, 0),
		(drawing, 313, 0, 4095, 0, 0),
		(drawing, 314, 0, 4095, 0, 0),
		(drawing, 315, 0, 4095, 0, 0),
		(drawing, 316, 0, 4095, 0, 0),
		(drawing, 317, 0, 4095, 0, 0),
		(drawing, 318, 0, 4095, 0, 0),
		(drawing, 319, 0, 4095, 0, 0),
		(drawing, 320, 0, 4095, 0, 0),
		(drawing, 321, 0, 4095, 0, 0),
		(drawing, 322, 0, 4095, 0, 0),
		(drawing, 323, 0, 4095, 0, 0),
		(drawing, 324, 0, 4095, 0, 0),
		(drawing, 325, 0, 4095, 0, 0),
		(drawing, 326, 0, 4095, 0, 0),
		(drawing, 327, 0, 4095, 0, 0),
		(drawing, 328, 0, 4095, 0, 0),
		(drawing, 329, 0, 4095, 0, 0),
		(drawing, 330, 0, 4095, 0, 0),
		(drawing, 331, 0, 4095, 0, 0),
		(drawing, 332, 0, 4095, 0, 0),
		(drawing, 333, 0, 4095, 0, 0),
		(drawing, 334, 0, 4095, 0, 0),
		(drawing, 335, 0, 4095, 0, 0),
		(drawing, 336, 0, 4095, 0, 0),
		(drawing, 337, 0, 4095, 0, 0),
		(drawing, 338, 0, 4095, 0, 0),
		(drawing, 339, 0, 4095, 0, 0),
		(drawing, 340, 0, 4095, 0, 0),
		(drawing, 341, 0, 4095, 0, 0),
		(drawing, 342, 0, 4095, 0, 0),
		(drawing, 343, 0, 4095, 0, 0),
		(drawing, 344, 0, 4095, 0, 0),
		(drawing, 345, 0, 4095, 0, 0),
		(drawing, 346, 0, 4095, 0, 0),
		(drawing, 347, 0, 4095, 0, 0),
		(drawing, 348, 0, 4095, 0, 0),
		(drawing, 349, 0, 4095, 0, 0),
		(drawing, 350, 0, 4095, 0, 0),
		(drawing, 351, 0, 4095, 0, 0),
		(drawing, 352, 0, 4095, 0, 0),
		(drawing, 353, 0, 4095, 0, 0),
		(drawing, 354, 0, 4095, 0, 0),
		(drawing, 355, 0, 4095, 0, 0),
		(drawing, 356, 0, 4095, 0, 0),
		(drawing, 357, 0, 4095, 0, 0),
		(drawing, 358, 0, 4095, 0, 0),
		(drawing, 359, 0, 4095, 0, 0),
		(drawing, 360, 0, 4095, 0, 0),
		(drawing, 361, 0, 4095, 0, 0),
		(drawing, 362, 0, 4095, 0, 0),
		(drawing, 363, 0, 4095, 0, 0),
		(drawing, 364, 0, 4095, 0, 0),
		(drawing, 365, 0, 4095, 0, 0),
		(drawing, 366, 0, 4095, 0, 0),
		(drawing, 367, 0, 4095, 0, 0),
		(drawing, 368, 0, 4095, 0, 0),
		(drawing, 369, 0, 4095, 0, 0),
		(drawing, 370, 0, 4095, 0, 0),
		(drawing, 371, 0, 4095, 0, 0),
		(drawing, 372, 0, 4095, 0, 0),
		(drawing, 373, 0, 4095, 0, 0),
		(drawing, 374, 0, 4095, 0, 0),
		(drawing, 375, 0, 4095, 0, 0),
		(drawing, 376, 0, 4095, 0, 0),
		(drawing, 377, 0, 4095, 0, 0),
		(drawing, 378, 0, 4095, 0, 0),
		(drawing, 379, 0, 4095, 0, 0),
		(drawing, 380, 0, 4095, 0, 0),
		(drawing, 381, 0, 4095, 0, 0),
		(drawing, 382, 0, 4095, 0, 0),
		(drawing, 383, 0, 4095, 0, 0),
		(drawing, 384, 0, 4095, 0, 0),
		(drawing, 385, 0, 4095, 0, 0),
		(drawing, 386, 0, 4095, 0, 0),
		(drawing, 387, 0, 4095, 0, 0),
		(drawing, 388, 0, 4095, 0, 0),
		(drawing, 389, 0, 4095, 0, 0),
		(drawing, 390, 0, 4095, 0, 0),
		(drawing, 391, 0, 4095, 0, 0),
		(drawing, 392, 0, 4095, 0, 0),
		(drawing, 393, 0, 4095, 0, 0),
		(drawing, 394, 0, 4095, 0, 0),
		(drawing, 395, 0, 4095, 0, 0),
		(drawing, 396, 0, 4095, 0, 0),
		(drawing, 397, 0, 4095, 0, 0),
		(drawing, 398, 0, 4095, 0, 0),
		(drawing, 399, 0, 4095, 0, 0),
		(drawing, 400, 0, 4095, 0, 0),
		(drawing, 401, 0, 4095, 0, 0),
		(drawing, 402, 0, 4095, 0, 0),
		(drawing, 403, 0, 4095, 0, 0),
		(drawing, 404, 0, 4095, 0, 0),
		(drawing, 405, 0, 4095, 0, 0),
		(drawing, 406, 0, 4095, 0, 0),
		(drawing, 407, 0, 4095, 0, 0),
		(drawing, 408, 0, 4095, 0, 0),
		(drawing, 409, 0, 4095, 0, 0),
		(drawing, 410, 0, 4095, 0, 0),
		(drawing, 411, 0, 4095, 0, 0),
		(drawing, 412, 0, 4095, 0, 0),
		(drawing, 413, 0, 4095, 0, 0),
		(drawing, 414, 0, 4095, 0, 0),
		(drawing, 415, 0, 4095, 0, 0),
		(drawing, 416, 0, 4095, 0, 0),
		(drawing, 417, 0, 4095, 0, 0),
		(drawing, 418, 0, 4095, 0, 0),
		(drawing, 419, 0, 4095, 0, 0),
		(drawing, 420, 0, 4095, 0, 0),
		(drawing, 421, 0, 4095, 0, 0),
		(drawing, 422, 0, 4095, 0, 0),
		(drawing, 423, 0, 4095, 0, 0),
		(drawing, 424, 0, 4095, 0, 0),
		(drawing, 425, 0, 4095, 0, 0),
		(drawing, 426, 0, 4095, 0, 0),
		(drawing, 427, 0, 4095, 0, 0),
		(drawing, 428, 0, 4095, 0, 0),
		(drawing, 429, 0, 4095, 0, 0),
		(drawing, 430, 0, 4095, 0, 0),
		(drawing, 431, 0, 4095, 0, 0),
		(drawing, 432, 0, 4095, 0, 0),
		(drawing, 433, 0, 4095, 0, 0),
		(drawing, 434, 0, 4095, 0, 0),
		(drawing, 435, 0, 4095, 0, 0),
		(drawing, 436, 0, 4095, 0, 0),
		(drawing, 437, 0, 4095, 0, 0),
		(drawing, 438, 0, 4095, 0, 0),
		(drawing, 439, 0, 4095, 0, 0),
		(drawing, 440, 0, 4095, 0, 0),
		(drawing, 441, 0, 4095, 0, 0),
		(drawing, 442, 0, 4095, 0, 0),
		(drawing, 443, 0, 4095, 0, 0),
		(drawing, 444, 0, 4095, 0, 0),
		(drawing, 445, 0, 4095, 0, 0),
		(drawing, 446, 0, 4095, 0, 0),
		(drawing, 447, 0, 4095, 0, 0),
		(drawing, 448, 0, 4095, 0, 0),
		(drawing, 449, 0, 4095, 0, 0),
		(drawing, 450, 0, 4095, 0, 0),
		(drawing, 451, 0, 4095, 0, 0),
		(drawing, 452, 0, 4095, 0, 0),
		(drawing, 453, 0, 4095, 0, 0),
		(drawing, 454, 0, 4095, 0, 0),
		(drawing, 455, 0, 4095, 0, 0),
		(drawing, 456, 0, 4095, 0, 0),
		(drawing, 457, 0, 4095, 0, 0),
		(drawing, 458, 0, 4095, 0, 0),
		(drawing, 459, 0, 4095, 0, 0),
		(drawing, 460, 0, 4095, 0, 0),
		(drawing, 461, 0, 4095, 0, 0),
		(drawing, 462, 0, 4095, 0, 0),
		(drawing, 463, 0, 4095, 0, 0),
		(drawing, 464, 0, 4095, 0, 0),
		(drawing, 465, 0, 4095, 0, 0),
		(drawing, 466, 0, 4095, 0, 0),
		(drawing, 467, 0, 4095, 0, 0),
		(drawing, 468, 0, 4095, 0, 0),
		(drawing, 469, 0, 4095, 0, 0),
		(drawing, 470, 0, 4095, 0, 0),
		(drawing, 471, 0, 4095, 0, 0),
		(drawing, 472, 0, 4095, 0, 0),
		(drawing, 473, 0, 4095, 0, 0),
		(drawing, 474, 0, 4095, 0, 0),
		(drawing, 475, 0, 4095, 0, 0),
		(drawing, 476, 0, 4095, 0, 0),
		(drawing, 477, 0, 4095, 0, 0),
		(drawing, 478, 0, 4095, 0, 0),
		(drawing, 479, 0, 4095, 0, 0),
		(drawing, 480, 0, 4095, 0, 0),
		(drawing, 481, 0, 4095, 0, 0),
		(drawing, 482, 0, 4095, 0, 0),
		(drawing, 483, 0, 4095, 0, 0),
		(drawing, 484, 0, 4095, 0, 0),
		(drawing, 485, 0, 4095, 0, 0),
		(drawing, 486, 0, 4095, 0, 0),
		(drawing, 487, 0, 4095, 0, 0),
		(drawing, 488, 0, 4095, 0, 0),
		(drawing, 489, 0, 4095, 0, 0),
		(drawing, 490, 0, 4095, 0, 0),
		(drawing, 491, 0, 4095, 0, 0),
		(drawing, 492, 0, 4095, 0, 0),
		(drawing, 493, 0, 4095, 0, 0),
		(drawing, 494, 0, 4095, 0, 0),
		(drawing, 495, 0, 4095, 0, 0),
		(drawing, 496, 0, 4095, 0, 0),
		(drawing, 497, 0, 4095, 0, 0),
		(drawing, 498, 0, 4095, 0, 0),
		(drawing, 499, 0, 4095, 0, 0),
		(drawing, 500, 0, 4095, 0, 0),
		(drawing, 501, 0, 4095, 0, 0),
		(drawing, 502, 0, 4095, 0, 0),
		(drawing, 503, 0, 4095, 0, 0),
		(drawing, 504, 0, 4095, 0, 0),
		(drawing, 505, 0, 4095, 0, 0),
		(drawing, 506, 0, 4095, 0, 0),
		(drawing, 507, 0, 4095, 0, 0),
		(drawing, 508, 0, 4095, 0, 0),
		(drawing, 509, 0, 4095, 0, 0),
		(drawing, 510, 0, 4095, 0, 0),
		(drawing, 511, 0, 4095, 0, 0),
		(drawing, 512, 0, 4095, 0, 0),
		(drawing, 513, 0, 4095, 0, 0),
		(drawing, 514, 0, 4095, 0, 0),
		(drawing, 515, 0, 4095, 0, 0),
		(drawing, 516, 0, 4095, 0, 0),
		(drawing, 517, 0, 4095, 0, 0),
		(drawing, 518, 0, 4095, 0, 0),
		(drawing, 519, 0, 4095, 0, 0),
		(drawing, 520, 0, 4095, 0, 0),
		(drawing, 521, 0, 4095, 0, 0),
		(drawing, 522, 0, 4095, 0, 0),
		(drawing, 523, 0, 4095, 0, 0),
		(drawing, 524, 0, 4095, 0, 0),
		(drawing, 525, 0, 4095, 0, 0),
		(drawing, 526, 0, 4095, 0, 0),
		(drawing, 527, 0, 4095, 0, 0),
		(drawing, 528, 0, 4095, 0, 0),
		(drawing, 529, 0, 4095, 0, 0),
		(drawing, 530, 0, 4095, 0, 0),
		(drawing, 531, 0, 4095, 0, 0),
		(drawing, 532, 0, 4095, 0, 0),
		(drawing, 533, 0, 4095, 0, 0),
		(drawing, 534, 0, 4095, 0, 0),
		(drawing, 535, 0, 4095, 0, 0),
		(drawing, 536, 0, 4095, 0, 0),
		(drawing, 537, 0, 4095, 0, 0),
		(drawing, 538, 0, 4095, 0, 0),
		(drawing, 539, 0, 4095, 0, 0),
		(drawing, 540, 0, 4095, 0, 0),
		(drawing, 541, 0, 4095, 0, 0),
		(drawing, 542, 0, 4095, 0, 0),
		(drawing, 543, 0, 4095, 0, 0),
		(drawing, 544, 0, 4095, 0, 0),
		(drawing, 545, 0, 4095, 0, 0),
		(drawing, 546, 0, 4095, 0, 0),
		(drawing, 547, 0, 4095, 0, 0),
		(drawing, 548, 0, 4095, 0, 0),
		(drawing, 549, 0, 4095, 0, 0),
		(drawing, 550, 0, 4095, 0, 0),
		(drawing, 551, 0, 4095, 0, 0),
		(drawing, 552, 0, 4095, 0, 0),
		(drawing, 553, 0, 4095, 0, 0),
		(drawing, 554, 0, 4095, 0, 0),
		(drawing, 555, 0, 4095, 0, 0),
		(drawing, 556, 0, 4095, 0, 0),
		(drawing, 557, 0, 4095, 0, 0),
		(drawing, 558, 0, 4095, 0, 0),
		(drawing, 559, 0, 4095, 0, 0),
		(drawing, 560, 0, 4095, 0, 0),
		(drawing, 561, 0, 4095, 0, 0),
		(drawing, 562, 0, 4095, 0, 0),
		(drawing, 563, 0, 4095, 0, 0),
		(drawing, 564, 0, 4095, 0, 0),
		(drawing, 565, 0, 4095, 0, 0),
		(drawing, 566, 0, 4095, 0, 0),
		(drawing, 567, 0, 4095, 0, 0),
		(drawing, 568, 0, 4095, 0, 0),
		(drawing, 569, 0, 4095, 0, 0),
		(drawing, 570, 0, 4095, 0, 0),
		(drawing, 571, 0, 4095, 0, 0),
		(drawing, 572, 0, 4095, 0, 0),
		(drawing, 573, 0, 4095, 0, 0),
		(drawing, 574, 0, 4095, 0, 0),
		(drawing, 575, 0, 4095, 0, 0),
		(drawing, 576, 0, 4095, 0, 0),
		(drawing, 577, 0, 4095, 0, 0),
		(drawing, 578, 0, 4095, 0, 0),
		(drawing, 579, 0, 4095, 0, 0),
		(drawing, 580, 0, 4095, 0, 0),
		(drawing, 581, 0, 4095, 0, 0),
		(drawing, 582, 0, 4095, 0, 0),
		(drawing, 583, 0, 4095, 0, 0),
		(drawing, 584, 0, 4095, 0, 0),
		(drawing, 585, 0, 4095, 0, 0),
		(drawing, 586, 0, 4095, 0, 0),
		(drawing, 587, 0, 4095, 0, 0),
		(drawing, 588, 0, 4095, 0, 0),
		(drawing, 589, 0, 4095, 0, 0),
		(drawing, 590, 0, 4095, 0, 0),
		(drawing, 591, 0, 4095, 0, 0),
		(drawing, 592, 0, 4095, 0, 0),
		(drawing, 593, 0, 4095, 0, 0),
		(drawing, 594, 0, 4095, 0, 0),
		(drawing, 595, 0, 4095, 0, 0),
		(drawing, 596, 0, 4095, 0, 0),
		(drawing, 597, 0, 4095, 0, 0),
		(drawing, 598, 0, 4095, 0, 0),
		(drawing, 599, 0, 4095, 0, 0),
		(drawing, 600, 0, 4095, 0, 0),
		(drawing, 601, 0, 4095, 0, 0),
		(drawing, 602, 0, 4095, 0, 0),
		(drawing, 603, 0, 4095, 0, 0),
		(drawing, 604, 0, 4095, 0, 0),
		(drawing, 605, 0, 4095, 0, 0),
		(drawing, 606, 0, 4095, 0, 0),
		(drawing, 607, 0, 4095, 0, 0),
		(drawing, 608, 0, 4095, 0, 0),
		(drawing, 609, 0, 4095, 0, 0),
		(drawing, 610, 0, 4095, 0, 0),
		(drawing, 611, 0, 4095, 0, 0),
		(drawing, 612, 0, 4095, 0, 0),
		(drawing, 613, 0, 4095, 0, 0),
		(drawing, 614, 0, 4095, 0, 0),
		(drawing, 615, 0, 4095, 0, 0),
		(drawing, 616, 0, 4095, 0, 0),
		(drawing, 617, 0, 4095, 0, 0),
		(drawing, 618, 0, 4095, 0, 0),
		(drawing, 619, 0, 4095, 0, 0),
		(drawing, 620, 0, 4095, 0, 0),
		(drawing, 621, 0, 4095, 0, 0),
		(drawing, 622, 0, 4095, 0, 0),
		(drawing, 623, 0, 4095, 0, 0),
		(drawing, 624, 0, 4095, 0, 0),
		(drawing, 625, 0, 4095, 0, 0),
		(drawing, 626, 0, 4095, 0, 0),
		(drawing, 627, 0, 4095, 0, 0),
		(drawing, 628, 0, 4095, 0, 0),
		(drawing, 629, 0, 4095, 0, 0),
		(drawing, 630, 0, 4095, 0, 0),
		(drawing, 631, 0, 4095, 0, 0),
		(drawing, 632, 0, 4095, 0, 0),
		(drawing, 633, 0, 4095, 0, 0),
		(drawing, 634, 0, 4095, 0, 0),
		(drawing, 635, 0, 4095, 0, 0),
		(drawing, 636, 0, 4095, 0, 0),
		(drawing, 637, 0, 4095, 0, 0),
		(drawing, 638, 0, 4095, 0, 0),
		(drawing, 639, 0, 4095, 0, 0),
		(drawing, 640, 0, 4095, 0, 0),
		(drawing, 641, 0, 4095, 0, 0),
		(drawing, 642, 0, 4095, 0, 0),
		(drawing, 643, 0, 4095, 0, 0),
		(drawing, 644, 0, 4095, 0, 0),
		(drawing, 645, 0, 4095, 0, 0),
		(drawing, 646, 0, 4095, 0, 0),
		(drawing, 647, 0, 4095, 0, 0),
		(drawing, 648, 0, 4095, 0, 0),
		(drawing, 649, 0, 4095, 0, 0),
		(drawing, 650, 0, 4095, 0, 0),
		(drawing, 651, 0, 4095, 0, 0),
		(drawing, 652, 0, 4095, 0, 0),
		(drawing, 653, 0, 4095, 0, 0),
		(drawing, 654, 0, 4095, 0, 0),
		(drawing, 655, 0, 4095, 0, 0),
		(drawing, 656, 0, 4095, 0, 0),
		(drawing, 657, 0, 4095, 0, 0),
		(drawing, 658, 0, 4095, 0, 0),
		(drawing, 659, 0, 4095, 0, 0),
		(drawing, 660, 0, 4095, 0, 0),
		(drawing, 661, 0, 4095, 0, 0),
		(drawing, 662, 0, 4095, 0, 0),
		(drawing, 663, 0, 4095, 0, 0),
		(drawing, 664, 0, 4095, 0, 0),
		(drawing, 665, 0, 4095, 0, 0),
		(drawing, 666, 0, 4095, 0, 0),
		(drawing, 667, 0, 4095, 0, 0),
		(drawing, 668, 0, 4095, 0, 0),
		(drawing, 669, 0, 4095, 0, 0),
		(drawing, 670, 0, 4095, 0, 0),
		(drawing, 671, 0, 4095, 0, 0),
		(drawing, 672, 0, 4095, 0, 0),
		(drawing, 673, 0, 4095, 0, 0),
		(drawing, 674, 0, 4095, 0, 0),
		(drawing, 675, 0, 4095, 0, 0),
		(drawing, 676, 0, 4095, 0, 0),
		(drawing, 677, 0, 4095, 0, 0),
		(drawing, 678, 0, 4095, 0, 0),
		(drawing, 679, 0, 4095, 0, 0),
		(drawing, 680, 0, 4095, 0, 0),
		(drawing, 681, 0, 4095, 0, 0),
		(drawing, 682, 0, 4095, 0, 0),
		(drawing, 683, 0, 4095, 0, 0),
		(drawing, 684, 0, 4095, 0, 0),
		(drawing, 685, 0, 4095, 0, 0),
		(drawing, 686, 0, 4095, 0, 0),
		(drawing, 687, 0, 4095, 0, 0),
		(drawing, 688, 0, 4095, 0, 0),
		(drawing, 689, 0, 4095, 0, 0),
		(drawing, 690, 0, 4095, 0, 0),
		(drawing, 691, 0, 4095, 0, 0),
		(drawing, 692, 0, 4095, 0, 0),
		(drawing, 693, 0, 4095, 0, 0),
		(drawing, 694, 0, 4095, 0, 0),
		(drawing, 695, 0, 4095, 0, 0),
		(drawing, 696, 0, 4095, 0, 0),
		(drawing, 697, 0, 4095, 0, 0),
		(drawing, 698, 0, 4095, 0, 0),
		(drawing, 699, 0, 4095, 0, 0),
		(drawing, 700, 0, 4095, 0, 0),
		(drawing, 701, 0, 4095, 0, 0),
		(drawing, 702, 0, 4095, 0, 0),
		(drawing, 703, 0, 4095, 0, 0),
		(drawing, 704, 0, 4095, 0, 0),
		(drawing, 705, 0, 4095, 0, 0),
		(drawing, 706, 0, 4095, 0, 0),
		(drawing, 707, 0, 4095, 0, 0),
		(drawing, 708, 0, 4095, 0, 0),
		(drawing, 709, 0, 4095, 0, 0),
		(drawing, 710, 0, 4095, 0, 0),
		(drawing, 711, 0, 4095, 0, 0),
		(drawing, 712, 0, 4095, 0, 0),
		(drawing, 713, 0, 4095, 0, 0),
		(drawing, 714, 0, 4095, 0, 0),
		(drawing, 715, 0, 4095, 0, 0),
		(drawing, 716, 0, 4095, 0, 0),
		(drawing, 717, 0, 4095, 0, 0),
		(drawing, 718, 0, 4095, 0, 0),
		(drawing, 719, 0, 4095, 0, 0),
		(drawing, 720, 0, 4095, 0, 0),
		(drawing, 721, 0, 4095, 0, 0),
		(drawing, 722, 0, 4095, 0, 0),
		(drawing, 723, 0, 4095, 0, 0),
		(drawing, 724, 0, 4095, 0, 0),
		(drawing, 725, 0, 4095, 0, 0),
		(drawing, 726, 0, 4095, 0, 0),
		(drawing, 727, 0, 4095, 0, 0),
		(drawing, 728, 0, 4095, 0, 0),
		(drawing, 729, 0, 4095, 0, 0),
		(drawing, 730, 0, 4095, 0, 0),
		(drawing, 731, 0, 4095, 0, 0),
		(drawing, 732, 0, 4095, 0, 0),
		(drawing, 733, 0, 4095, 0, 0),
		(drawing, 734, 0, 4095, 0, 0),
		(drawing, 735, 0, 4095, 0, 0),
		(drawing, 736, 0, 4095, 0, 0),
		(drawing, 737, 0, 4095, 0, 0),
		(drawing, 738, 0, 4095, 0, 0),
		(drawing, 739, 0, 4095, 0, 0),
		(drawing, 740, 0, 4095, 0, 0),
		(drawing, 741, 0, 4095, 0, 0),
		(drawing, 742, 0, 4095, 0, 0),
		(drawing, 743, 0, 4095, 0, 0),
		(drawing, 744, 0, 4095, 0, 0),
		(drawing, 745, 0, 4095, 0, 0),
		(drawing, 746, 0, 4095, 0, 0),
		(drawing, 747, 0, 4095, 0, 0),
		(drawing, 748, 0, 4095, 0, 0),
		(drawing, 749, 0, 4095, 0, 0),
		(drawing, 750, 0, 4095, 0, 0),
		(drawing, 751, 0, 4095, 0, 0),
		(drawing, 752, 0, 4095, 0, 0),
		(drawing, 753, 0, 4095, 0, 0),
		(drawing, 754, 0, 4095, 0, 0),
		(drawing, 755, 0, 4095, 0, 0),
		(drawing, 756, 0, 4095, 0, 0),
		(drawing, 757, 0, 4095, 0, 0),
		(drawing, 758, 0, 4095, 0, 0),
		(drawing, 759, 0, 4095, 0, 0),
		(drawing, 760, 0, 4095, 0, 0),
		(drawing, 761, 0, 4095, 0, 0),
		(drawing, 762, 0, 4095, 0, 0),
		(drawing, 763, 0, 4095, 0, 0),
		(drawing, 764, 0, 4095, 0, 0),
		(drawing, 765, 0, 4095, 0, 0),
		(drawing, 766, 0, 4095, 0, 0),
		(drawing, 767, 0, 4095, 0, 0),
		(drawing, 768, 0, 4095, 0, 0),
		(drawing, 769, 0, 4095, 0, 0),
		(drawing, 770, 0, 4095, 0, 0),
		(drawing, 771, 0, 4095, 0, 0),
		(drawing, 772, 0, 4095, 0, 0),
		(drawing, 773, 0, 4095, 0, 0),
		(drawing, 774, 0, 4095, 0, 0),
		(drawing, 775, 0, 4095, 0, 0),
		(drawing, 776, 0, 4095, 0, 0),
		(drawing, 777, 0, 4095, 0, 0),
		(drawing, 778, 0, 4095, 0, 0),
		(drawing, 779, 0, 4095, 0, 0),
		(drawing, 780, 0, 4095, 0, 0),
		(drawing, 781, 0, 4095, 0, 0),
		(drawing, 782, 0, 4095, 0, 0),
		(drawing, 783, 0, 4095, 0, 0),
		(drawing, 784, 0, 4095, 0, 0),
		(drawing, 785, 0, 4095, 0, 0),
		(drawing, 786, 0, 4095, 0, 0),
		(drawing, 787, 0, 4095, 0, 0),
		(drawing, 788, 0, 4095, 0, 0),
		(drawing, 789, 0, 4095, 0, 0),
		(drawing, 790, 0, 4095, 0, 0),
		(drawing, 791, 0, 4095, 0, 0),
		(drawing, 792, 0, 4095, 0, 0),
		(drawing, 793, 0, 4095, 0, 0),
		(drawing, 794, 0, 4095, 0, 0),
		(drawing, 795, 0, 4095, 0, 0),
		(drawing, 796, 0, 4095, 0, 0),
		(drawing, 797, 0, 4095, 0, 0),
		(drawing, 798, 0, 4095, 0, 0),
		(drawing, 799, 0, 4095, 0, 0),
		(drawing, 800, 0, 4095, 0, 0),
		(drawing, 801, 0, 4095, 0, 0),
		(drawing, 802, 0, 4095, 0, 0),
		(drawing, 803, 0, 4095, 0, 0),
		(drawing, 804, 0, 4095, 0, 0),
		(drawing, 805, 0, 4095, 0, 0),
		(drawing, 806, 0, 4095, 0, 0),
		(drawing, 807, 0, 4095, 0, 0),
		(drawing, 808, 0, 4095, 0, 0),
		(drawing, 809, 0, 4095, 0, 0),
		(drawing, 810, 0, 4095, 0, 0),
		(drawing, 811, 0, 4095, 0, 0),
		(drawing, 812, 0, 4095, 0, 0),
		(drawing, 813, 0, 4095, 0, 0),
		(drawing, 814, 0, 4095, 0, 0),
		(drawing, 815, 0, 4095, 0, 0),
		(drawing, 816, 0, 4095, 0, 0),
		(drawing, 817, 0, 4095, 0, 0),
		(drawing, 818, 0, 4095, 0, 0),
		(drawing, 819, 0, 4095, 0, 0),
		(drawing, 820, 0, 4095, 0, 0),
		(drawing, 821, 0, 4095, 0, 0),
		(drawing, 822, 0, 4095, 0, 0),
		(drawing, 823, 0, 4095, 0, 0),
		(drawing, 824, 0, 4095, 0, 0),
		(drawing, 825, 0, 4095, 0, 0),
		(drawing, 826, 0, 4095, 0, 0),
		(drawing, 827, 0, 4095, 0, 0),
		(drawing, 828, 0, 4095, 0, 0),
		(drawing, 829, 0, 4095, 0, 0),
		(drawing, 830, 0, 4095, 0, 0),
		(drawing, 831, 0, 4095, 0, 0),
		(drawing, 832, 0, 4095, 0, 0),
		(drawing, 833, 0, 4095, 0, 0),
		(drawing, 834, 0, 4095, 0, 0),
		(drawing, 835, 0, 4095, 0, 0),
		(drawing, 836, 0, 4095, 0, 0),
		(drawing, 837, 0, 4095, 0, 0),
		(drawing, 838, 0, 4095, 0, 0),
		(drawing, 839, 0, 4095, 0, 0),
		(drawing, 840, 0, 4095, 0, 0),
		(drawing, 841, 0, 4095, 0, 0),
		(drawing, 842, 0, 4095, 0, 0),
		(drawing, 843, 0, 4095, 0, 0),
		(drawing, 844, 0, 4095, 0, 0),
		(drawing, 845, 0, 4095, 0, 0),
		(drawing, 846, 0, 4095, 0, 0),
		(drawing, 847, 0, 4095, 0, 0),
		(drawing, 848, 0, 4095, 0, 0),
		(drawing, 849, 0, 4095, 0, 0),
		(drawing, 850, 0, 4095, 0, 0),
		(drawing, 851, 0, 4095, 0, 0),
		(drawing, 852, 0, 4095, 0, 0),
		(drawing, 853, 0, 4095, 0, 0),
		(drawing, 854, 0, 4095, 0, 0),
		(drawing, 855, 0, 4095, 0, 0),
		(drawing, 856, 0, 4095, 0, 0),
		(drawing, 857, 0, 4095, 0, 0),
		(drawing, 858, 0, 4095, 0, 0),
		(drawing, 859, 0, 4095, 0, 0),
		(drawing, 860, 0, 4095, 0, 0),
		(drawing, 861, 0, 4095, 0, 0),
		(drawing, 862, 0, 4095, 0, 0),
		(drawing, 863, 0, 4095, 0, 0),
		(drawing, 864, 0, 4095, 0, 0),
		(drawing, 865, 0, 4095, 0, 0),
		(drawing, 866, 0, 4095, 0, 0),
		(drawing, 867, 0, 4095, 0, 0),
		(drawing, 868, 0, 4095, 0, 0),
		(drawing, 869, 0, 4095, 0, 0),
		(drawing, 870, 0, 4095, 0, 0),
		(drawing, 871, 0, 4095, 0, 0),
		(drawing, 872, 0, 4095, 0, 0),
		(drawing, 873, 0, 4095, 0, 0),
		(drawing, 874, 0, 4095, 0, 0),
		(drawing, 875, 0, 4095, 0, 0),
		(drawing, 876, 0, 4095, 0, 0),
		(drawing, 877, 0, 4095, 0, 0),
		(drawing, 878, 0, 4095, 0, 0),
		(drawing, 879, 0, 4095, 0, 0),
		(drawing, 880, 0, 4095, 0, 0),
		(drawing, 881, 0, 4095, 0, 0),
		(drawing, 882, 0, 4095, 0, 0),
		(drawing, 883, 0, 4095, 0, 0),
		(drawing, 884, 0, 4095, 0, 0),
		(drawing, 885, 0, 4095, 0, 0),
		(drawing, 886, 0, 4095, 0, 0),
		(drawing, 887, 0, 4095, 0, 0),
		(drawing, 888, 0, 4095, 0, 0),
		(drawing, 889, 0, 4095, 0, 0),
		(drawing, 890, 0, 4095, 0, 0),
		(drawing, 891, 0, 4095, 0, 0),
		(drawing, 892, 0, 4095, 0, 0),
		(drawing, 893, 0, 4095, 0, 0),
		(drawing, 894, 0, 4095, 0, 0),
		(drawing, 895, 0, 4095, 0, 0),
		(drawing, 896, 0, 4095, 0, 0),
		(drawing, 897, 0, 4095, 0, 0),
		(drawing, 898, 0, 4095, 0, 0),
		(drawing, 899, 0, 4095, 0, 0),
		(drawing, 900, 0, 4095, 0, 0),
		(drawing, 901, 0, 4095, 0, 0),
		(drawing, 902, 0, 4095, 0, 0),
		(drawing, 903, 0, 4095, 0, 0),
		(drawing, 904, 0, 4095, 0, 0),
		(drawing, 905, 0, 4095, 0, 0),
		(drawing, 906, 0, 4095, 0, 0),
		(drawing, 907, 0, 4095, 0, 0),
		(drawing, 908, 0, 4095, 0, 0),
		(drawing, 909, 0, 4095, 0, 0),
		(drawing, 910, 0, 4095, 0, 0),
		(drawing, 911, 0, 4095, 0, 0),
		(drawing, 912, 0, 4095, 0, 0),
		(drawing, 913, 0, 4095, 0, 0),
		(drawing, 914, 0, 4095, 0, 0),
		(drawing, 915, 0, 4095, 0, 0),
		(drawing, 916, 0, 4095, 0, 0),
		(drawing, 917, 0, 4095, 0, 0),
		(drawing, 918, 0, 4095, 0, 0),
		(drawing, 919, 0, 4095, 0, 0),
		(drawing, 920, 0, 4095, 0, 0),
		(drawing, 921, 0, 4095, 0, 0),
		(drawing, 922, 0, 4095, 0, 0),
		(drawing, 923, 0, 4095, 0, 0),
		(drawing, 924, 0, 4095, 0, 0),
		(drawing, 925, 0, 4095, 0, 0),
		(drawing, 926, 0, 4095, 0, 0),
		(drawing, 927, 0, 4095, 0, 0),
		(drawing, 928, 0, 4095, 0, 0),
		(drawing, 929, 0, 4095, 0, 0),
		(drawing, 930, 0, 4095, 0, 0),
		(drawing, 931, 0, 4095, 0, 0),
		(drawing, 932, 0, 4095, 0, 0),
		(drawing, 933, 0, 4095, 0, 0),
		(drawing, 934, 0, 4095, 0, 0),
		(drawing, 935, 0, 4095, 0, 0),
		(drawing, 936, 0, 4095, 0, 0),
		(drawing, 937, 0, 4095, 0, 0),
		(drawing, 938, 0, 4095, 0, 0),
		(drawing, 939, 0, 4095, 0, 0),
		(drawing, 940, 0, 4095, 0, 0),
		(drawing, 941, 0, 4095, 0, 0),
		(drawing, 942, 0, 4095, 0, 0),
		(drawing, 943, 0, 4095, 0, 0),
		(drawing, 944, 0, 4095, 0, 0),
		(drawing, 945, 0, 4095, 0, 0),
		(drawing, 946, 0, 4095, 0, 0),
		(drawing, 947, 0, 4095, 0, 0),
		(drawing, 948, 0, 4095, 0, 0),
		(drawing, 949, 0, 4095, 0, 0),
		(drawing, 950, 0, 4095, 0, 0),
		(drawing, 951, 0, 4095, 0, 0),
		(drawing, 952, 0, 4095, 0, 0),
		(drawing, 953, 0, 4095, 0, 0),
		(drawing, 954, 0, 4095, 0, 0),
		(drawing, 955, 0, 4095, 0, 0),
		(drawing, 956, 0, 4095, 0, 0),
		(drawing, 957, 0, 4095, 0, 0),
		(drawing, 958, 0, 4095, 0, 0),
		(drawing, 959, 0, 4095, 0, 0),
		(drawing, 960, 0, 4095, 0, 0),
		(drawing, 961, 0, 4095, 0, 0),
		(drawing, 962, 0, 4095, 0, 0),
		(drawing, 963, 0, 4095, 0, 0),
		(drawing, 964, 0, 4095, 0, 0),
		(drawing, 965, 0, 4095, 0, 0),
		(drawing, 966, 0, 4095, 0, 0),
		(drawing, 967, 0, 4095, 0, 0),
		(drawing, 968, 0, 4095, 0, 0),
		(drawing, 969, 0, 4095, 0, 0),
		(drawing, 970, 0, 4095, 0, 0),
		(drawing, 971, 0, 4095, 0, 0),
		(drawing, 972, 0, 4095, 0, 0),
		(drawing, 973, 0, 4095, 0, 0),
		(drawing, 974, 0, 4095, 0, 0),
		(drawing, 975, 0, 4095, 0, 0),
		(drawing, 976, 0, 4095, 0, 0),
		(drawing, 977, 0, 4095, 0, 0),
		(drawing, 978, 0, 4095, 0, 0),
		(drawing, 979, 0, 4095, 0, 0),
		(drawing, 980, 0, 4095, 0, 0),
		(drawing, 981, 0, 4095, 0, 0),
		(drawing, 982, 0, 4095, 0, 0),
		(drawing, 983, 0, 4095, 0, 0),
		(drawing, 984, 0, 4095, 0, 0),
		(drawing, 985, 0, 4095, 0, 0),
		(drawing, 986, 0, 4095, 0, 0),
		(drawing, 987, 0, 4095, 0, 0),
		(drawing, 988, 0, 4095, 0, 0),
		(drawing, 989, 0, 4095, 0, 0),
		(drawing, 990, 0, 4095, 0, 0),
		(drawing, 991, 0, 4095, 0, 0),
		(drawing, 992, 0, 4095, 0, 0),
		(drawing, 993, 0, 4095, 0, 0),
		(drawing, 994, 0, 4095, 0, 0),
		(drawing, 995, 0, 4095, 0, 0),
		(drawing, 996, 0, 4095, 0, 0),
		(drawing, 997, 0, 4095, 0, 0),
		(drawing, 998, 0, 4095, 0, 0),
		(drawing, 999, 0, 4095, 0, 0),
		(drawing, 1000, 0, 4095, 0, 0),
		(drawing, 1001, 0, 4095, 0, 0),
		(drawing, 1002, 0, 4095, 0, 0),
		(drawing, 1003, 0, 4095, 0, 0),
		(drawing, 1004, 0, 4095, 0, 0),
		(drawing, 1005, 0, 4095, 0, 0),
		(drawing, 1006, 0, 4095, 0, 0),
		(drawing, 1007, 0, 4095, 0, 0),
		(drawing, 1008, 0, 4095, 0, 0),
		(drawing, 1009, 0, 4095, 0, 0),
		(drawing, 1010, 0, 4095, 0, 0),
		(drawing, 1011, 0, 4095, 0, 0),
		(drawing, 1012, 0, 4095, 0, 0),
		(drawing, 1013, 0, 4095, 0, 0),
		(drawing, 1014, 0, 4095, 0, 0),
		(drawing, 1015, 0, 4095, 0, 0),
		(drawing, 1016, 0, 4095, 0, 0),
		(drawing, 1017, 0, 4095, 0, 0),
		(drawing, 1018, 0, 4095, 0, 0),
		(drawing, 1019, 0, 4095, 0, 0),
		(drawing, 1020, 0, 4095, 0, 0),
		(drawing, 1021, 0, 4095, 0, 0),
		(drawing, 1022, 0, 4095, 0, 0),
		(drawing, 1023, 0, 4095, 0, 0),
		(drawing, 1024, 0, 4095, 0, 0),
		(drawing, 1025, 0, 4095, 0, 0),
		(drawing, 1026, 0, 4095, 0, 0),
		(drawing, 1027, 0, 4095, 0, 0),
		(drawing, 1028, 0, 4095, 0, 0),
		(drawing, 1029, 0, 4095, 0, 0),
		(drawing, 1030, 0, 4095, 0, 0),
		(drawing, 1031, 0, 4095, 0, 0),
		(drawing, 1032, 0, 4095, 0, 0),
		(drawing, 1033, 0, 4095, 0, 0),
		(drawing, 1034, 0, 4095, 0, 0),
		(drawing, 1035, 0, 4095, 0, 0),
		(drawing, 1036, 0, 4095, 0, 0),
		(drawing, 1037, 0, 4095, 0, 0),
		(drawing, 1038, 0, 4095, 0, 0),
		(drawing, 1039, 0, 4095, 0, 0),
		(drawing, 1040, 0, 4095, 0, 0),
		(drawing, 1041, 0, 4095, 0, 0),
		(drawing, 1042, 0, 4095, 0, 0),
		(drawing, 1043, 0, 4095, 0, 0),
		(drawing, 1044, 0, 4095, 0, 0),
		(drawing, 1045, 0, 4095, 0, 0),
		(drawing, 1046, 0, 4095, 0, 0),
		(drawing, 1047, 0, 4095, 0, 0),
		(drawing, 1048, 0, 4095, 0, 0),
		(drawing, 1049, 0, 4095, 0, 0),
		(drawing, 1050, 0, 4095, 0, 0),
		(drawing, 1051, 0, 4095, 0, 0),
		(drawing, 1052, 0, 4095, 0, 0),
		(drawing, 1053, 0, 4095, 0, 0),
		(drawing, 1054, 0, 4095, 0, 0),
		(drawing, 1055, 0, 4095, 0, 0),
		(drawing, 1056, 0, 4095, 0, 0),
		(drawing, 1057, 0, 4095, 0, 0),
		(drawing, 1058, 0, 4095, 0, 0),
		(drawing, 1059, 0, 4095, 0, 0),
		(drawing, 1060, 0, 4095, 0, 0),
		(drawing, 1061, 0, 4095, 0, 0),
		(drawing, 1062, 0, 4095, 0, 0),
		(drawing, 1063, 0, 4095, 0, 0),
		(drawing, 1064, 0, 4095, 0, 0),
		(drawing, 1065, 0, 4095, 0, 0),
		(drawing, 1066, 0, 4095, 0, 0),
		(drawing, 1067, 0, 4095, 0, 0),
		(drawing, 1068, 0, 4095, 0, 0),
		(drawing, 1069, 0, 4095, 0, 0),
		(drawing, 1070, 0, 4095, 0, 0),
		(drawing, 1071, 0, 4095, 0, 0),
		(drawing, 1072, 0, 4095, 0, 0),
		(drawing, 1073, 0, 4095, 0, 0),
		(drawing, 1074, 0, 4095, 0, 0),
		(drawing, 1075, 0, 4095, 0, 0),
		(drawing, 1076, 0, 4095, 0, 0),
		(drawing, 1077, 0, 4095, 0, 0),
		(drawing, 1078, 0, 4095, 0, 0),
		(drawing, 1079, 0, 4095, 0, 0),
		(drawing, 1080, 0, 4095, 0, 0),
		(drawing, 1081, 0, 4095, 0, 0),
		(drawing, 1082, 0, 4095, 0, 0),
		(drawing, 1083, 0, 4095, 0, 0),
		(drawing, 1084, 0, 4095, 0, 0),
		(drawing, 1085, 0, 4095, 0, 0),
		(drawing, 1086, 0, 4095, 0, 0),
		(drawing, 1087, 0, 4095, 0, 0),
		(drawing, 1088, 0, 4095, 0, 0),
		(drawing, 1089, 0, 4095, 0, 0),
		(drawing, 1090, 0, 4095, 0, 0),
		(drawing, 1091, 0, 4095, 0, 0),
		(drawing, 1092, 0, 4095, 0, 0),
		(drawing, 1093, 0, 4095, 0, 0),
		(drawing, 1094, 0, 4095, 0, 0),
		(drawing, 1095, 0, 4095, 0, 0),
		(drawing, 1096, 0, 4095, 0, 0),
		(drawing, 1097, 0, 4095, 0, 0),
		(drawing, 1098, 0, 4095, 0, 0),
		(drawing, 1099, 0, 4095, 0, 0),
		(drawing, 1100, 0, 4095, 0, 0),
		(drawing, 1101, 0, 4095, 0, 0),
		(drawing, 1102, 0, 4095, 0, 0),
		(drawing, 1103, 0, 4095, 0, 0),
		(drawing, 1104, 0, 4095, 0, 0),
		(drawing, 1105, 0, 4095, 0, 0),
		(drawing, 1106, 0, 4095, 0, 0),
		(drawing, 1107, 0, 4095, 0, 0),
		(drawing, 1108, 0, 4095, 0, 0),
		(drawing, 1109, 0, 4095, 0, 0),
		(drawing, 1110, 0, 4095, 0, 0),
		(drawing, 1111, 0, 4095, 0, 0),
		(drawing, 1112, 0, 4095, 0, 0),
		(drawing, 1113, 0, 4095, 0, 0),
		(drawing, 1114, 0, 4095, 0, 0),
		(drawing, 1115, 0, 4095, 0, 0),
		(drawing, 1116, 0, 4095, 0, 0),
		(drawing, 1117, 0, 4095, 0, 0),
		(drawing, 1118, 0, 4095, 0, 0),
		(drawing, 1119, 0, 4095, 0, 0),
		(drawing, 1120, 0, 4095, 0, 0),
		(drawing, 1121, 0, 4095, 0, 0),
		(drawing, 1122, 0, 4095, 0, 0),
		(drawing, 1123, 0, 4095, 0, 0),
		(drawing, 1124, 0, 4095, 0, 0),
		(drawing, 1125, 0, 4095, 0, 0),
		(drawing, 1126, 0, 4095, 0, 0),
		(drawing, 1127, 0, 4095, 0, 0),
		(drawing, 1128, 0, 4095, 0, 0),
		(drawing, 1129, 0, 4095, 0, 0),
		(drawing, 1130, 0, 4095, 0, 0),
		(drawing, 1131, 0, 4095, 0, 0),
		(drawing, 1132, 0, 4095, 0, 0),
		(drawing, 1133, 0, 4095, 0, 0),
		(drawing, 1134, 0, 4095, 0, 0),
		(drawing, 1135, 0, 4095, 0, 0),
		(drawing, 1136, 0, 4095, 0, 0),
		(drawing, 1137, 0, 4095, 0, 0),
		(drawing, 1138, 0, 4095, 0, 0),
		(drawing, 1139, 0, 4095, 0, 0),
		(drawing, 1140, 0, 4095, 0, 0),
		(drawing, 1141, 0, 4095, 0, 0),
		(drawing, 1142, 0, 4095, 0, 0),
		(drawing, 1143, 0, 4095, 0, 0),
		(drawing, 1144, 0, 4095, 0, 0),
		(drawing, 1145, 0, 4095, 0, 0),
		(drawing, 1146, 0, 4095, 0, 0),
		(drawing, 1147, 0, 4095, 0, 0),
		(drawing, 1148, 0, 4095, 0, 0),
		(drawing, 1149, 0, 4095, 0, 0),
		(drawing, 1150, 0, 4095, 0, 0),
		(drawing, 1151, 0, 4095, 0, 0),
		(drawing, 1152, 0, 4095, 0, 0),
		(drawing, 1153, 0, 4095, 0, 0),
		(drawing, 1154, 0, 4095, 0, 0),
		(drawing, 1155, 0, 4095, 0, 0),
		(drawing, 1156, 0, 4095, 0, 0),
		(drawing, 1157, 0, 4095, 0, 0),
		(drawing, 1158, 0, 4095, 0, 0),
		(drawing, 1159, 0, 4095, 0, 0),
		(drawing, 1160, 0, 4095, 0, 0),
		(drawing, 1161, 0, 4095, 0, 0),
		(drawing, 1162, 0, 4095, 0, 0),
		(drawing, 1163, 0, 4095, 0, 0),
		(drawing, 1164, 0, 4095, 0, 0),
		(drawing, 1165, 0, 4095, 0, 0),
		(drawing, 1166, 0, 4095, 0, 0),
		(drawing, 1167, 0, 4095, 0, 0),
		(drawing, 1168, 0, 4095, 0, 0),
		(drawing, 1169, 0, 4095, 0, 0),
		(drawing, 1170, 0, 4095, 0, 0),
		(drawing, 1171, 0, 4095, 0, 0),
		(drawing, 1172, 0, 4095, 0, 0),
		(drawing, 1173, 0, 4095, 0, 0),
		(drawing, 1174, 0, 4095, 0, 0),
		(drawing, 1175, 0, 4095, 0, 0),
		(drawing, 1176, 0, 4095, 0, 0),
		(drawing, 1177, 0, 4095, 0, 0),
		(drawing, 1178, 0, 4095, 0, 0),
		(drawing, 1179, 0, 4095, 0, 0),
		(drawing, 1180, 0, 4095, 0, 0),
		(drawing, 1181, 0, 4095, 0, 0),
		(drawing, 1182, 0, 4095, 0, 0),
		(drawing, 1183, 0, 4095, 0, 0),
		(drawing, 1184, 0, 4095, 0, 0),
		(drawing, 1185, 0, 4095, 0, 0),
		(drawing, 1186, 0, 4095, 0, 0),
		(drawing, 1187, 0, 4095, 0, 0),
		(drawing, 1188, 0, 4095, 0, 0),
		(drawing, 1189, 0, 4095, 0, 0),
		(drawing, 1190, 0, 4095, 0, 0),
		(drawing, 1191, 0, 4095, 0, 0),
		(drawing, 1192, 0, 4095, 0, 0),
		(drawing, 1193, 0, 4095, 0, 0),
		(drawing, 1194, 0, 4095, 0, 0),
		(drawing, 1195, 0, 4095, 0, 0),
		(drawing, 1196, 0, 4095, 0, 0),
		(drawing, 1197, 0, 4095, 0, 0),
		(drawing, 1198, 0, 4095, 0, 0),
		(drawing, 1199, 0, 4095, 0, 0),
		(drawing, 1200, 0, 4095, 0, 0),
		(drawing, 1201, 0, 4095, 0, 0),
		(drawing, 1202, 0, 4095, 0, 0),
		(drawing, 1203, 0, 4095, 0, 0),
		(drawing, 1204, 0, 4095, 0, 0),
		(drawing, 1205, 0, 4095, 0, 0),
		(drawing, 1206, 0, 4095, 0, 0),
		(drawing, 1207, 0, 4095, 0, 0),
		(drawing, 1208, 0, 4095, 0, 0),
		(drawing, 1209, 0, 4095, 0, 0),
		(drawing, 1210, 0, 4095, 0, 0),
		(drawing, 1211, 0, 4095, 0, 0),
		(drawing, 1212, 0, 4095, 0, 0),
		(drawing, 1213, 0, 4095, 0, 0),
		(drawing, 1214, 0, 4095, 0, 0),
		(drawing, 1215, 0, 4095, 0, 0),
		(drawing, 1216, 0, 4095, 0, 0),
		(drawing, 1217, 0, 4095, 0, 0),
		(drawing, 1218, 0, 4095, 0, 0),
		(drawing, 1219, 0, 4095, 0, 0),
		(drawing, 1220, 0, 4095, 0, 0),
		(drawing, 1221, 0, 4095, 0, 0),
		(drawing, 1222, 0, 4095, 0, 0),
		(drawing, 1223, 0, 4095, 0, 0),
		(drawing, 1224, 0, 4095, 0, 0),
		(drawing, 1225, 0, 4095, 0, 0),
		(drawing, 1226, 0, 4095, 0, 0),
		(drawing, 1227, 0, 4095, 0, 0),
		(drawing, 1228, 0, 4095, 0, 0),
		(drawing, 1229, 0, 4095, 0, 0),
		(drawing, 1230, 0, 4095, 0, 0),
		(drawing, 1231, 0, 4095, 0, 0),
		(drawing, 1232, 0, 4095, 0, 0),
		(drawing, 1233, 0, 4095, 0, 0),
		(drawing, 1234, 0, 4095, 0, 0),
		(drawing, 1235, 0, 4095, 0, 0),
		(drawing, 1236, 0, 4095, 0, 0),
		(drawing, 1237, 0, 4095, 0, 0),
		(drawing, 1238, 0, 4095, 0, 0),
		(drawing, 1239, 0, 4095, 0, 0),
		(drawing, 1240, 0, 4095, 0, 0),
		(drawing, 1241, 0, 4095, 0, 0),
		(drawing, 1242, 0, 4095, 0, 0),
		(drawing, 1243, 0, 4095, 0, 0),
		(drawing, 1244, 0, 4095, 0, 0),
		(drawing, 1245, 0, 4095, 0, 0),
		(drawing, 1246, 0, 4095, 0, 0),
		(drawing, 1247, 0, 4095, 0, 0),
		(drawing, 1248, 0, 4095, 0, 0),
		(drawing, 1249, 0, 4095, 0, 0),
		(drawing, 1250, 0, 4095, 0, 0),
		(drawing, 1251, 0, 4095, 0, 0),
		(drawing, 1252, 0, 4095, 0, 0),
		(drawing, 1253, 0, 4095, 0, 0),
		(drawing, 1254, 0, 4095, 0, 0),
		(drawing, 1255, 0, 4095, 0, 0),
		(drawing, 1256, 0, 4095, 0, 0),
		(drawing, 1257, 0, 4095, 0, 0),
		(drawing, 1258, 0, 4095, 0, 0),
		(drawing, 1259, 0, 4095, 0, 0),
		(drawing, 1260, 0, 4095, 0, 0),
		(drawing, 1261, 0, 4095, 0, 0),
		(drawing, 1262, 0, 4095, 0, 0),
		(drawing, 1263, 0, 4095, 0, 0),
		(drawing, 1264, 0, 4095, 0, 0),
		(drawing, 1265, 0, 4095, 0, 0),
		(drawing, 1266, 0, 4095, 0, 0),
		(drawing, 1267, 0, 4095, 0, 0),
		(drawing, 1268, 0, 4095, 0, 0),
		(drawing, 1269, 0, 4095, 0, 0),
		(drawing, 1270, 0, 4095, 0, 0),
		(drawing, 1271, 0, 4095, 0, 0),
		(drawing, 1272, 0, 4095, 0, 0),
		(drawing, 1273, 0, 4095, 0, 0),
		(drawing, 1274, 0, 4095, 0, 0),
		(drawing, 1275, 0, 4095, 0, 0),
		(drawing, 1276, 0, 4095, 0, 0),
		(drawing, 1277, 0, 4095, 0, 0),
		(drawing, 1278, 0, 4095, 0, 0),
		(drawing, 1279, 0, 4095, 0, 0),
		(drawing, 1280, 0, 4095, 0, 0),
		(drawing, 1281, 0, 4095, 0, 0),
		(drawing, 1282, 0, 4095, 0, 0),
		(drawing, 1283, 0, 4095, 0, 0),
		(drawing, 1284, 0, 4095, 0, 0),
		(drawing, 1285, 0, 4095, 0, 0),
		(drawing, 1286, 0, 4095, 0, 0),
		(drawing, 1287, 0, 4095, 0, 0),
		(drawing, 1288, 0, 4095, 0, 0),
		(drawing, 1289, 0, 4095, 0, 0),
		(drawing, 1290, 0, 4095, 0, 0),
		(drawing, 1291, 0, 4095, 0, 0),
		(drawing, 1292, 0, 4095, 0, 0),
		(drawing, 1293, 0, 4095, 0, 0),
		(drawing, 1294, 0, 4095, 0, 0),
		(drawing, 1295, 0, 4095, 0, 0),
		(drawing, 1296, 0, 4095, 0, 0),
		(drawing, 1297, 0, 4095, 0, 0),
		(drawing, 1298, 0, 4095, 0, 0),
		(drawing, 1299, 0, 4095, 0, 0),
		(drawing, 1300, 0, 4095, 0, 0),
		(drawing, 1301, 0, 4095, 0, 0),
		(drawing, 1302, 0, 4095, 0, 0),
		(drawing, 1303, 0, 4095, 0, 0),
		(drawing, 1304, 0, 4095, 0, 0),
		(drawing, 1305, 0, 4095, 0, 0),
		(drawing, 1306, 0, 4095, 0, 0),
		(drawing, 1307, 0, 4095, 0, 0),
		(drawing, 1308, 0, 4095, 0, 0),
		(drawing, 1309, 0, 4095, 0, 0),
		(drawing, 1310, 0, 4095, 0, 0),
		(drawing, 1311, 0, 4095, 0, 0),
		(drawing, 1312, 0, 4095, 0, 0),
		(drawing, 1313, 0, 4095, 0, 0),
		(drawing, 1314, 0, 4095, 0, 0),
		(drawing, 1315, 0, 4095, 0, 0),
		(drawing, 1316, 0, 4095, 0, 0),
		(drawing, 1317, 0, 4095, 0, 0),
		(drawing, 1318, 0, 4095, 0, 0),
		(drawing, 1319, 0, 4095, 0, 0),
		(drawing, 1320, 0, 4095, 0, 0),
		(drawing, 1321, 0, 4095, 0, 0),
		(drawing, 1322, 0, 4095, 0, 0),
		(drawing, 1323, 0, 4095, 0, 0),
		(drawing, 1324, 0, 4095, 0, 0),
		(drawing, 1325, 0, 4095, 0, 0),
		(drawing, 1326, 0, 4095, 0, 0),
		(drawing, 1327, 0, 4095, 0, 0),
		(drawing, 1328, 0, 4095, 0, 0),
		(drawing, 1329, 0, 4095, 0, 0),
		(drawing, 1330, 0, 4095, 0, 0),
		(drawing, 1331, 0, 4095, 0, 0),
		(drawing, 1332, 0, 4095, 0, 0),
		(drawing, 1333, 0, 4095, 0, 0),
		(drawing, 1334, 0, 4095, 0, 0),
		(drawing, 1335, 0, 4095, 0, 0),
		(drawing, 1336, 0, 4095, 0, 0),
		(drawing, 1337, 0, 4095, 0, 0),
		(drawing, 1338, 0, 4095, 0, 0),
		(drawing, 1339, 0, 4095, 0, 0),
		(drawing, 1340, 0, 4095, 0, 0),
		(drawing, 1341, 0, 4095, 0, 0),
		(drawing, 1342, 0, 4095, 0, 0),
		(drawing, 1343, 0, 4095, 0, 0),
		(drawing, 1344, 0, 4095, 0, 0),
		(drawing, 1345, 0, 4095, 0, 0),
		(drawing, 1346, 0, 4095, 0, 0),
		(drawing, 1347, 0, 4095, 0, 0),
		(drawing, 1348, 0, 4095, 0, 0),
		(drawing, 1349, 0, 4095, 0, 0),
		(drawing, 1350, 0, 4095, 0, 0),
		(drawing, 1351, 0, 4095, 0, 0),
		(drawing, 1352, 0, 4095, 0, 0),
		(drawing, 1353, 0, 4095, 0, 0),
		(drawing, 1354, 0, 4095, 0, 0),
		(drawing, 1355, 0, 4095, 0, 0),
		(drawing, 1356, 0, 4095, 0, 0),
		(drawing, 1357, 0, 4095, 0, 0),
		(drawing, 1358, 0, 4095, 0, 0),
		(drawing, 1359, 0, 4095, 0, 0),
		(drawing, 1360, 0, 4095, 0, 0),
		(drawing, 1361, 0, 4095, 0, 0),
		(drawing, 1362, 0, 4095, 0, 0),
		(drawing, 1363, 0, 4095, 0, 0),
		(drawing, 1364, 0, 4095, 0, 0),
		(drawing, 1365, 0, 4095, 0, 0),
		(drawing, 1366, 0, 4095, 0, 0),
		(drawing, 1367, 0, 4095, 0, 0),
		(drawing, 1368, 0, 4095, 0, 0),
		(drawing, 1369, 0, 4095, 0, 0),
		(drawing, 1370, 0, 4095, 0, 0),
		(drawing, 1371, 0, 4095, 0, 0),
		(drawing, 1372, 0, 4095, 0, 0),
		(drawing, 1373, 0, 4095, 0, 0),
		(drawing, 1374, 0, 4095, 0, 0),
		(drawing, 1375, 0, 4095, 0, 0),
		(drawing, 1376, 0, 4095, 0, 0),
		(drawing, 1377, 0, 4095, 0, 0),
		(drawing, 1378, 0, 4095, 0, 0),
		(drawing, 1379, 0, 4095, 0, 0),
		(drawing, 1380, 0, 4095, 0, 0),
		(drawing, 1381, 0, 4095, 0, 0),
		(drawing, 1382, 0, 4095, 0, 0),
		(drawing, 1383, 0, 4095, 0, 0),
		(drawing, 1384, 0, 4095, 0, 0),
		(drawing, 1385, 0, 4095, 0, 0),
		(drawing, 1386, 0, 4095, 0, 0),
		(drawing, 1387, 0, 4095, 0, 0),
		(drawing, 1388, 0, 4095, 0, 0),
		(drawing, 1389, 0, 4095, 0, 0),
		(drawing, 1390, 0, 4095, 0, 0),
		(drawing, 1391, 0, 4095, 0, 0),
		(drawing, 1392, 0, 4095, 0, 0),
		(drawing, 1393, 0, 4095, 0, 0),
		(drawing, 1394, 0, 4095, 0, 0),
		(drawing, 1395, 0, 4095, 0, 0),
		(drawing, 1396, 0, 4095, 0, 0),
		(drawing, 1397, 0, 4095, 0, 0),
		(drawing, 1398, 0, 4095, 0, 0),
		(drawing, 1399, 0, 4095, 0, 0),
		(drawing, 1400, 0, 4095, 0, 0),
		(drawing, 1401, 0, 4095, 0, 0),
		(drawing, 1402, 0, 4095, 0, 0),
		(drawing, 1403, 0, 4095, 0, 0),
		(drawing, 1404, 0, 4095, 0, 0),
		(drawing, 1405, 0, 4095, 0, 0),
		(drawing, 1406, 0, 4095, 0, 0),
		(drawing, 1407, 0, 4095, 0, 0),
		(drawing, 1408, 0, 4095, 0, 0),
		(drawing, 1409, 0, 4095, 0, 0),
		(drawing, 1410, 0, 4095, 0, 0),
		(drawing, 1411, 0, 4095, 0, 0),
		(drawing, 1412, 0, 4095, 0, 0),
		(drawing, 1413, 0, 4095, 0, 0),
		(drawing, 1414, 0, 4095, 0, 0),
		(drawing, 1415, 0, 4095, 0, 0),
		(drawing, 1416, 0, 4095, 0, 0),
		(drawing, 1417, 0, 4095, 0, 0),
		(drawing, 1418, 0, 4095, 0, 0),
		(drawing, 1419, 0, 4095, 0, 0),
		(drawing, 1420, 0, 4095, 0, 0),
		(drawing, 1421, 0, 4095, 0, 0),
		(drawing, 1422, 0, 4095, 0, 0),
		(drawing, 1423, 0, 4095, 0, 0),
		(drawing, 1424, 0, 4095, 0, 0),
		(drawing, 1425, 0, 4095, 0, 0),
		(drawing, 1426, 0, 4095, 0, 0),
		(drawing, 1427, 0, 4095, 0, 0),
		(drawing, 1428, 0, 4095, 0, 0),
		(drawing, 1429, 0, 4095, 0, 0),
		(drawing, 1430, 0, 4095, 0, 0),
		(drawing, 1431, 0, 4095, 0, 0),
		(drawing, 1432, 0, 4095, 0, 0),
		(drawing, 1433, 0, 4095, 0, 0),
		(drawing, 1434, 0, 4095, 0, 0),
		(drawing, 1435, 0, 4095, 0, 0),
		(drawing, 1436, 0, 4095, 0, 0),
		(drawing, 1437, 0, 4095, 0, 0),
		(drawing, 1438, 0, 4095, 0, 0),
		(drawing, 1439, 0, 4095, 0, 0),
		(drawing, 1440, 0, 4095, 0, 0),
		(drawing, 1441, 0, 4095, 0, 0),
		(drawing, 1442, 0, 4095, 0, 0),
		(drawing, 1443, 0, 4095, 0, 0),
		(drawing, 1444, 0, 4095, 0, 0),
		(drawing, 1445, 0, 4095, 0, 0),
		(drawing, 1446, 0, 4095, 0, 0),
		(drawing, 1447, 0, 4095, 0, 0),
		(drawing, 1448, 0, 4095, 0, 0),
		(drawing, 1449, 0, 4095, 0, 0),
		(drawing, 1450, 0, 4095, 0, 0),
		(drawing, 1451, 0, 4095, 0, 0),
		(drawing, 1452, 0, 4095, 0, 0),
		(drawing, 1453, 0, 4095, 0, 0),
		(drawing, 1454, 0, 4095, 0, 0),
		(drawing, 1455, 0, 4095, 0, 0),
		(drawing, 1456, 0, 4095, 0, 0),
		(drawing, 1457, 0, 4095, 0, 0),
		(drawing, 1458, 0, 4095, 0, 0),
		(drawing, 1459, 0, 4095, 0, 0),
		(drawing, 1460, 0, 4095, 0, 0),
		(drawing, 1461, 0, 4095, 0, 0),
		(drawing, 1462, 0, 4095, 0, 0),
		(drawing, 1463, 0, 4095, 0, 0),
		(drawing, 1464, 0, 4095, 0, 0),
		(drawing, 1465, 0, 4095, 0, 0),
		(drawing, 1466, 0, 4095, 0, 0),
		(drawing, 1467, 0, 4095, 0, 0),
		(drawing, 1468, 0, 4095, 0, 0),
		(drawing, 1469, 0, 4095, 0, 0),
		(drawing, 1470, 0, 4095, 0, 0),
		(drawing, 1471, 0, 4095, 0, 0),
		(drawing, 1472, 0, 4095, 0, 0),
		(drawing, 1473, 0, 4095, 0, 0),
		(drawing, 1474, 0, 4095, 0, 0),
		(drawing, 1475, 0, 4095, 0, 0),
		(drawing, 1476, 0, 4095, 0, 0),
		(drawing, 1477, 0, 4095, 0, 0),
		(drawing, 1478, 0, 4095, 0, 0),
		(drawing, 1479, 0, 4095, 0, 0),
		(drawing, 1480, 0, 4095, 0, 0),
		(drawing, 1481, 0, 4095, 0, 0),
		(drawing, 1482, 0, 4095, 0, 0),
		(drawing, 1483, 0, 4095, 0, 0),
		(drawing, 1484, 0, 4095, 0, 0),
		(drawing, 1485, 0, 4095, 0, 0),
		(drawing, 1486, 0, 4095, 0, 0),
		(drawing, 1487, 0, 4095, 0, 0),
		(drawing, 1488, 0, 4095, 0, 0),
		(drawing, 1489, 0, 4095, 0, 0),
		(drawing, 1490, 0, 4095, 0, 0),
		(drawing, 1491, 0, 4095, 0, 0),
		(drawing, 1492, 0, 4095, 0, 0),
		(drawing, 1493, 0, 4095, 0, 0),
		(drawing, 1494, 0, 4095, 0, 0),
		(drawing, 1495, 0, 4095, 0, 0),
		(drawing, 1496, 0, 4095, 0, 0),
		(drawing, 1497, 0, 4095, 0, 0),
		(drawing, 1498, 0, 4095, 0, 0),
		(drawing, 1499, 0, 4095, 0, 0),
		(drawing, 1500, 0, 4095, 0, 0),
		(drawing, 1501, 0, 4095, 0, 0),
		(drawing, 1502, 0, 4095, 0, 0),
		(drawing, 1503, 0, 4095, 0, 0),
		(drawing, 1504, 0, 4095, 0, 0),
		(drawing, 1505, 0, 4095, 0, 0),
		(drawing, 1506, 0, 4095, 0, 0),
		(drawing, 1507, 0, 4095, 0, 0),
		(drawing, 1508, 0, 4095, 0, 0),
		(drawing, 1509, 0, 4095, 0, 0),
		(drawing, 1510, 0, 4095, 0, 0),
		(drawing, 1511, 0, 4095, 0, 0),
		(drawing, 1512, 0, 4095, 0, 0),
		(drawing, 1513, 0, 4095, 0, 0),
		(drawing, 1514, 0, 4095, 0, 0),
		(drawing, 1515, 0, 4095, 0, 0),
		(drawing, 1516, 0, 4095, 0, 0),
		(drawing, 1517, 0, 4095, 0, 0),
		(drawing, 1518, 0, 4095, 0, 0),
		(drawing, 1519, 0, 4095, 0, 0),
		(drawing, 1520, 0, 4095, 0, 0),
		(drawing, 1521, 0, 4095, 0, 0),
		(drawing, 1522, 0, 4095, 0, 0),
		(drawing, 1523, 0, 4095, 0, 0),
		(drawing, 1524, 0, 4095, 0, 0),
		(drawing, 1525, 0, 4095, 0, 0),
		(drawing, 1526, 0, 4095, 0, 0),
		(drawing, 1527, 0, 4095, 0, 0),
		(drawing, 1528, 0, 4095, 0, 0),
		(drawing, 1529, 0, 4095, 0, 0),
		(drawing, 1530, 0, 4095, 0, 0),
		(drawing, 1531, 0, 4095, 0, 0),
		(drawing, 1532, 0, 4095, 0, 0),
		(drawing, 1533, 0, 4095, 0, 0),
		(drawing, 1534, 0, 4095, 0, 0),
		(drawing, 1535, 0, 4095, 0, 0),
		(drawing, 1536, 0, 4095, 0, 0),
		(drawing, 1537, 0, 4095, 0, 0),
		(drawing, 1538, 0, 4095, 0, 0),
		(drawing, 1539, 0, 4095, 0, 0),
		(drawing, 1540, 0, 4095, 0, 0),
		(drawing, 1541, 0, 4095, 0, 0),
		(drawing, 1542, 0, 4095, 0, 0),
		(drawing, 1543, 0, 4095, 0, 0),
		(drawing, 1544, 0, 4095, 0, 0),
		(drawing, 1545, 0, 4095, 0, 0),
		(drawing, 1546, 0, 4095, 0, 0),
		(drawing, 1547, 0, 4095, 0, 0),
		(drawing, 1548, 0, 4095, 0, 0),
		(drawing, 1549, 0, 4095, 0, 0),
		(drawing, 1550, 0, 4095, 0, 0),
		(drawing, 1551, 0, 4095, 0, 0),
		(drawing, 1552, 0, 4095, 0, 0),
		(drawing, 1553, 0, 4095, 0, 0),
		(drawing, 1554, 0, 4095, 0, 0),
		(drawing, 1555, 0, 4095, 0, 0),
		(drawing, 1556, 0, 4095, 0, 0),
		(drawing, 1557, 0, 4095, 0, 0),
		(drawing, 1558, 0, 4095, 0, 0),
		(drawing, 1559, 0, 4095, 0, 0),
		(drawing, 1560, 0, 4095, 0, 0),
		(drawing, 1561, 0, 4095, 0, 0),
		(drawing, 1562, 0, 4095, 0, 0),
		(drawing, 1563, 0, 4095, 0, 0),
		(drawing, 1564, 0, 4095, 0, 0),
		(drawing, 1565, 0, 4095, 0, 0),
		(drawing, 1566, 0, 4095, 0, 0),
		(drawing, 1567, 0, 4095, 0, 0),
		(drawing, 1568, 0, 4095, 0, 0),
		(drawing, 1569, 0, 4095, 0, 0),
		(drawing, 1570, 0, 4095, 0, 0),
		(drawing, 1571, 0, 4095, 0, 0),
		(drawing, 1572, 0, 4095, 0, 0),
		(drawing, 1573, 0, 4095, 0, 0),
		(drawing, 1574, 0, 4095, 0, 0),
		(drawing, 1575, 0, 4095, 0, 0),
		(drawing, 1576, 0, 4095, 0, 0),
		(drawing, 1577, 0, 4095, 0, 0),
		(drawing, 1578, 0, 4095, 0, 0),
		(drawing, 1579, 0, 4095, 0, 0),
		(drawing, 1580, 0, 4095, 0, 0),
		(drawing, 1581, 0, 4095, 0, 0),
		(drawing, 1582, 0, 4095, 0, 0),
		(drawing, 1583, 0, 4095, 0, 0),
		(drawing, 1584, 0, 4095, 0, 0),
		(drawing, 1585, 0, 4095, 0, 0),
		(drawing, 1586, 0, 4095, 0, 0),
		(drawing, 1587, 0, 4095, 0, 0),
		(drawing, 1588, 0, 4095, 0, 0),
		(drawing, 1589, 0, 4095, 0, 0),
		(drawing, 1590, 0, 4095, 0, 0),
		(drawing, 1591, 0, 4095, 0, 0),
		(drawing, 1592, 0, 4095, 0, 0),
		(drawing, 1593, 0, 4095, 0, 0),
		(drawing, 1594, 0, 4095, 0, 0),
		(drawing, 1595, 0, 4095, 0, 0),
		(drawing, 1596, 0, 4095, 0, 0),
		(drawing, 1597, 0, 4095, 0, 0),
		(drawing, 1598, 0, 4095, 0, 0),
		(drawing, 1599, 0, 4095, 0, 0),
		(drawing, 1600, 0, 4095, 0, 0),
		(drawing, 1601, 0, 4095, 0, 0),
		(drawing, 1602, 0, 4095, 0, 0),
		(drawing, 1603, 0, 4095, 0, 0),
		(drawing, 1604, 0, 4095, 0, 0),
		(drawing, 1605, 0, 4095, 0, 0),
		(drawing, 1606, 0, 4095, 0, 0),
		(drawing, 1607, 0, 4095, 0, 0),
		(drawing, 1608, 0, 4095, 0, 0),
		(drawing, 1609, 0, 4095, 0, 0),
		(drawing, 1610, 0, 4095, 0, 0),
		(drawing, 1611, 0, 4095, 0, 0),
		(drawing, 1612, 0, 4095, 0, 0),
		(drawing, 1613, 0, 4095, 0, 0),
		(drawing, 1614, 0, 4095, 0, 0),
		(drawing, 1615, 0, 4095, 0, 0),
		(drawing, 1616, 0, 4095, 0, 0),
		(drawing, 1617, 0, 4095, 0, 0),
		(drawing, 1618, 0, 4095, 0, 0),
		(drawing, 1619, 0, 4095, 0, 0),
		(drawing, 1620, 0, 4095, 0, 0),
		(drawing, 1621, 0, 4095, 0, 0),
		(drawing, 1622, 0, 4095, 0, 0),
		(drawing, 1623, 0, 4095, 0, 0),
		(drawing, 1624, 0, 4095, 0, 0),
		(drawing, 1625, 0, 4095, 0, 0),
		(drawing, 1626, 0, 4095, 0, 0),
		(drawing, 1627, 0, 4095, 0, 0),
		(drawing, 1628, 0, 4095, 0, 0),
		(drawing, 1629, 0, 4095, 0, 0),
		(drawing, 1630, 0, 4095, 0, 0),
		(drawing, 1631, 0, 4095, 0, 0),
		(drawing, 1632, 0, 4095, 0, 0),
		(drawing, 1633, 0, 4095, 0, 0),
		(drawing, 1634, 0, 4095, 0, 0),
		(drawing, 1635, 0, 4095, 0, 0),
		(drawing, 1636, 0, 4095, 0, 0),
		(drawing, 1637, 0, 4095, 0, 0),
		(drawing, 1638, 0, 4095, 0, 0),
		(drawing, 1639, 0, 4095, 0, 0),
		(drawing, 1640, 0, 4095, 0, 0),
		(drawing, 1641, 0, 4095, 0, 0),
		(drawing, 1642, 0, 4095, 0, 0),
		(drawing, 1643, 0, 4095, 0, 0),
		(drawing, 1644, 0, 4095, 0, 0),
		(drawing, 1645, 0, 4095, 0, 0),
		(drawing, 1646, 0, 4095, 0, 0),
		(drawing, 1647, 0, 4095, 0, 0),
		(drawing, 1648, 0, 4095, 0, 0),
		(drawing, 1649, 0, 4095, 0, 0),
		(drawing, 1650, 0, 4095, 0, 0),
		(drawing, 1651, 0, 4095, 0, 0),
		(drawing, 1652, 0, 4095, 0, 0),
		(drawing, 1653, 0, 4095, 0, 0),
		(drawing, 1654, 0, 4095, 0, 0),
		(drawing, 1655, 0, 4095, 0, 0),
		(drawing, 1656, 0, 4095, 0, 0),
		(drawing, 1657, 0, 4095, 0, 0),
		(drawing, 1658, 0, 4095, 0, 0),
		(drawing, 1659, 0, 4095, 0, 0),
		(drawing, 1660, 0, 4095, 0, 0),
		(drawing, 1661, 0, 4095, 0, 0),
		(drawing, 1662, 0, 4095, 0, 0),
		(drawing, 1663, 0, 4095, 0, 0),
		(drawing, 1664, 0, 4095, 0, 0),
		(drawing, 1665, 0, 4095, 0, 0),
		(drawing, 1666, 0, 4095, 0, 0),
		(drawing, 1667, 0, 4095, 0, 0),
		(drawing, 1668, 0, 4095, 0, 0),
		(drawing, 1669, 0, 4095, 0, 0),
		(drawing, 1670, 0, 4095, 0, 0),
		(drawing, 1671, 0, 4095, 0, 0),
		(drawing, 1672, 0, 4095, 0, 0),
		(drawing, 1673, 0, 4095, 0, 0),
		(drawing, 1674, 0, 4095, 0, 0),
		(drawing, 1675, 0, 4095, 0, 0),
		(drawing, 1676, 0, 4095, 0, 0),
		(drawing, 1677, 0, 4095, 0, 0),
		(drawing, 1678, 0, 4095, 0, 0),
		(drawing, 1679, 0, 4095, 0, 0),
		(drawing, 1680, 0, 4095, 0, 0),
		(drawing, 1681, 0, 4095, 0, 0),
		(drawing, 1682, 0, 4095, 0, 0),
		(drawing, 1683, 0, 4095, 0, 0),
		(drawing, 1684, 0, 4095, 0, 0),
		(drawing, 1685, 0, 4095, 0, 0),
		(drawing, 1686, 0, 4095, 0, 0),
		(drawing, 1687, 0, 4095, 0, 0),
		(drawing, 1688, 0, 4095, 0, 0),
		(drawing, 1689, 0, 4095, 0, 0),
		(drawing, 1690, 0, 4095, 0, 0),
		(drawing, 1691, 0, 4095, 0, 0),
		(drawing, 1692, 0, 4095, 0, 0),
		(drawing, 1693, 0, 4095, 0, 0),
		(drawing, 1694, 0, 4095, 0, 0),
		(drawing, 1695, 0, 4095, 0, 0),
		(drawing, 1696, 0, 4095, 0, 0),
		(drawing, 1697, 0, 4095, 0, 0),
		(drawing, 1698, 0, 4095, 0, 0),
		(drawing, 1699, 0, 4095, 0, 0),
		(drawing, 1700, 0, 4095, 0, 0),
		(drawing, 1701, 0, 4095, 0, 0),
		(drawing, 1702, 0, 4095, 0, 0),
		(drawing, 1703, 0, 4095, 0, 0),
		(drawing, 1704, 0, 4095, 0, 0),
		(drawing, 1705, 0, 4095, 0, 0),
		(drawing, 1706, 0, 4095, 0, 0),
		(drawing, 1707, 0, 4095, 0, 0),
		(drawing, 1708, 0, 4095, 0, 0),
		(drawing, 1709, 0, 4095, 0, 0),
		(drawing, 1710, 0, 4095, 0, 0),
		(drawing, 1711, 0, 4095, 0, 0),
		(drawing, 1712, 0, 4095, 0, 0),
		(drawing, 1713, 0, 4095, 0, 0),
		(drawing, 1714, 0, 4095, 0, 0),
		(drawing, 1715, 0, 4095, 0, 0),
		(drawing, 1716, 0, 4095, 0, 0),
		(drawing, 1717, 0, 4095, 0, 0),
		(drawing, 1718, 0, 4095, 0, 0),
		(drawing, 1719, 0, 4095, 0, 0),
		(drawing, 1720, 0, 4095, 0, 0),
		(drawing, 1721, 0, 4095, 0, 0),
		(drawing, 1722, 0, 4095, 0, 0),
		(drawing, 1723, 0, 4095, 0, 0),
		(drawing, 1724, 0, 4095, 0, 0),
		(drawing, 1725, 0, 4095, 0, 0),
		(drawing, 1726, 0, 4095, 0, 0),
		(drawing, 1727, 0, 4095, 0, 0),
		(drawing, 1728, 0, 4095, 0, 0),
		(drawing, 1729, 0, 4095, 0, 0),
		(drawing, 1730, 0, 4095, 0, 0),
		(drawing, 1731, 0, 4095, 0, 0),
		(drawing, 1732, 0, 4095, 0, 0),
		(drawing, 1733, 0, 4095, 0, 0),
		(drawing, 1734, 0, 4095, 0, 0),
		(drawing, 1735, 0, 4095, 0, 0),
		(drawing, 1736, 0, 4095, 0, 0),
		(drawing, 1737, 0, 4095, 0, 0),
		(drawing, 1738, 0, 4095, 0, 0),
		(drawing, 1739, 0, 4095, 0, 0),
		(drawing, 1740, 0, 4095, 0, 0),
		(drawing, 1741, 0, 4095, 0, 0),
		(drawing, 1742, 0, 4095, 0, 0),
		(drawing, 1743, 0, 4095, 0, 0),
		(drawing, 1744, 0, 4095, 0, 0),
		(drawing, 1745, 0, 4095, 0, 0),
		(drawing, 1746, 0, 4095, 0, 0),
		(drawing, 1747, 0, 4095, 0, 0),
		(drawing, 1748, 0, 4095, 0, 0),
		(drawing, 1749, 0, 4095, 0, 0),
		(drawing, 1750, 0, 4095, 0, 0),
		(drawing, 1751, 0, 4095, 0, 0),
		(drawing, 1752, 0, 4095, 0, 0),
		(drawing, 1753, 0, 4095, 0, 0),
		(drawing, 1754, 0, 4095, 0, 0),
		(drawing, 1755, 0, 4095, 0, 0),
		(drawing, 1756, 0, 4095, 0, 0),
		(drawing, 1757, 0, 4095, 0, 0),
		(drawing, 1758, 0, 4095, 0, 0),
		(drawing, 1759, 0, 4095, 0, 0),
		(drawing, 1760, 0, 4095, 0, 0),
		(drawing, 1761, 0, 4095, 0, 0),
		(drawing, 1762, 0, 4095, 0, 0),
		(drawing, 1763, 0, 4095, 0, 0),
		(drawing, 1764, 0, 4095, 0, 0),
		(drawing, 1765, 0, 4095, 0, 0),
		(drawing, 1766, 0, 4095, 0, 0),
		(drawing, 1767, 0, 4095, 0, 0),
		(drawing, 1768, 0, 4095, 0, 0),
		(drawing, 1769, 0, 4095, 0, 0),
		(drawing, 1770, 0, 4095, 0, 0),
		(drawing, 1771, 0, 4095, 0, 0),
		(drawing, 1772, 0, 4095, 0, 0),
		(drawing, 1773, 0, 4095, 0, 0),
		(drawing, 1774, 0, 4095, 0, 0),
		(drawing, 1775, 0, 4095, 0, 0),
		(drawing, 1776, 0, 4095, 0, 0),
		(drawing, 1777, 0, 4095, 0, 0),
		(drawing, 1778, 0, 4095, 0, 0),
		(drawing, 1779, 0, 4095, 0, 0),
		(drawing, 1780, 0, 4095, 0, 0),
		(drawing, 1781, 0, 4095, 0, 0),
		(drawing, 1782, 0, 4095, 0, 0),
		(drawing, 1783, 0, 4095, 0, 0),
		(drawing, 1784, 0, 4095, 0, 0),
		(drawing, 1785, 0, 4095, 0, 0),
		(drawing, 1786, 0, 4095, 0, 0),
		(drawing, 1787, 0, 4095, 0, 0),
		(drawing, 1788, 0, 4095, 0, 0),
		(drawing, 1789, 0, 4095, 0, 0),
		(drawing, 1790, 0, 4095, 0, 0),
		(drawing, 1791, 0, 4095, 0, 0),
		(drawing, 1792, 0, 4095, 0, 0),
		(drawing, 1793, 0, 4095, 0, 0),
		(drawing, 1794, 0, 4095, 0, 0),
		(drawing, 1795, 0, 4095, 0, 0),
		(drawing, 1796, 0, 4095, 0, 0),
		(drawing, 1797, 0, 4095, 0, 0),
		(drawing, 1798, 0, 4095, 0, 0),
		(drawing, 1799, 0, 4095, 0, 0),
		(drawing, 1800, 0, 4095, 0, 0),
		(drawing, 1801, 0, 4095, 0, 0),
		(drawing, 1802, 0, 4095, 0, 0),
		(drawing, 1803, 0, 4095, 0, 0),
		(drawing, 1804, 0, 4095, 0, 0),
		(drawing, 1805, 0, 4095, 0, 0),
		(drawing, 1806, 0, 4095, 0, 0),
		(drawing, 1807, 0, 4095, 0, 0),
		(drawing, 1808, 0, 4095, 0, 0),
		(drawing, 1809, 0, 4095, 0, 0),
		(drawing, 1810, 0, 4095, 0, 0),
		(drawing, 1811, 0, 4095, 0, 0),
		(drawing, 1812, 0, 4095, 0, 0),
		(drawing, 1813, 0, 4095, 0, 0),
		(drawing, 1814, 0, 4095, 0, 0),
		(drawing, 1815, 0, 4095, 0, 0),
		(drawing, 1816, 0, 4095, 0, 0),
		(drawing, 1817, 0, 4095, 0, 0),
		(drawing, 1818, 0, 4095, 0, 0),
		(drawing, 1819, 0, 4095, 0, 0),
		(drawing, 1820, 0, 4095, 0, 0),
		(drawing, 1821, 0, 4095, 0, 0),
		(drawing, 1822, 0, 4095, 0, 0),
		(drawing, 1823, 0, 4095, 0, 0),
		(drawing, 1824, 0, 4095, 0, 0),
		(drawing, 1825, 0, 4095, 0, 0),
		(drawing, 1826, 0, 4095, 0, 0),
		(drawing, 1827, 0, 4095, 0, 0),
		(drawing, 1828, 0, 4095, 0, 0),
		(drawing, 1829, 0, 4095, 0, 0),
		(drawing, 1830, 0, 4095, 0, 0),
		(drawing, 1831, 0, 4095, 0, 0),
		(drawing, 1832, 0, 4095, 0, 0),
		(drawing, 1833, 0, 4095, 0, 0),
		(drawing, 1834, 0, 4095, 0, 0),
		(drawing, 1835, 0, 4095, 0, 0),
		(drawing, 1836, 0, 4095, 0, 0),
		(drawing, 1837, 0, 4095, 0, 0),
		(drawing, 1838, 0, 4095, 0, 0),
		(drawing, 1839, 0, 4095, 0, 0),
		(drawing, 1840, 0, 4095, 0, 0),
		(drawing, 1841, 0, 4095, 0, 0),
		(drawing, 1842, 0, 4095, 0, 0),
		(drawing, 1843, 0, 4095, 0, 0),
		(drawing, 1844, 0, 4095, 0, 0),
		(drawing, 1845, 0, 4095, 0, 0),
		(drawing, 1846, 0, 4095, 0, 0),
		(drawing, 1847, 0, 4095, 0, 0),
		(drawing, 1848, 0, 4095, 0, 0),
		(drawing, 1849, 0, 4095, 0, 0),
		(drawing, 1850, 0, 4095, 0, 0),
		(drawing, 1851, 0, 4095, 0, 0),
		(drawing, 1852, 0, 4095, 0, 0),
		(drawing, 1853, 0, 4095, 0, 0),
		(drawing, 1854, 0, 4095, 0, 0),
		(drawing, 1855, 0, 4095, 0, 0),
		(drawing, 1856, 0, 4095, 0, 0),
		(drawing, 1857, 0, 4095, 0, 0),
		(drawing, 1858, 0, 4095, 0, 0),
		(drawing, 1859, 0, 4095, 0, 0),
		(drawing, 1860, 0, 4095, 0, 0),
		(drawing, 1861, 0, 4095, 0, 0),
		(drawing, 1862, 0, 4095, 0, 0),
		(drawing, 1863, 0, 4095, 0, 0),
		(drawing, 1864, 0, 4095, 0, 0),
		(drawing, 1865, 0, 4095, 0, 0),
		(drawing, 1866, 0, 4095, 0, 0),
		(drawing, 1867, 0, 4095, 0, 0),
		(drawing, 1868, 0, 4095, 0, 0),
		(drawing, 1869, 0, 4095, 0, 0),
		(drawing, 1870, 0, 4095, 0, 0),
		(drawing, 1871, 0, 4095, 0, 0),
		(drawing, 1872, 0, 4095, 0, 0),
		(drawing, 1873, 0, 4095, 0, 0),
		(drawing, 1874, 0, 4095, 0, 0),
		(drawing, 1875, 0, 4095, 0, 0),
		(drawing, 1876, 0, 4095, 0, 0),
		(drawing, 1877, 0, 4095, 0, 0),
		(drawing, 1878, 0, 4095, 0, 0),
		(drawing, 1879, 0, 4095, 0, 0),
		(drawing, 1880, 0, 4095, 0, 0),
		(drawing, 1881, 0, 4095, 0, 0),
		(drawing, 1882, 0, 4095, 0, 0),
		(drawing, 1883, 0, 4095, 0, 0),
		(drawing, 1884, 0, 4095, 0, 0),
		(drawing, 1885, 0, 4095, 0, 0),
		(drawing, 1886, 0, 4095, 0, 0),
		(drawing, 1887, 0, 4095, 0, 0),
		(drawing, 1888, 0, 4095, 0, 0),
		(drawing, 1889, 0, 4095, 0, 0),
		(drawing, 1890, 0, 4095, 0, 0),
		(drawing, 1891, 0, 4095, 0, 0),
		(drawing, 1892, 0, 4095, 0, 0),
		(drawing, 1893, 0, 4095, 0, 0),
		(drawing, 1894, 0, 4095, 0, 0),
		(drawing, 1895, 0, 4095, 0, 0),
		(drawing, 1896, 0, 4095, 0, 0),
		(drawing, 1897, 0, 4095, 0, 0),
		(drawing, 1898, 0, 4095, 0, 0),
		(drawing, 1899, 0, 4095, 0, 0),
		(drawing, 1900, 0, 4095, 0, 0),
		(drawing, 1901, 0, 4095, 0, 0),
		(drawing, 1902, 0, 4095, 0, 0),
		(drawing, 1903, 0, 4095, 0, 0),
		(drawing, 1904, 0, 4095, 0, 0),
		(drawing, 1905, 0, 4095, 0, 0),
		(drawing, 1906, 0, 4095, 0, 0),
		(drawing, 1907, 0, 4095, 0, 0),
		(drawing, 1908, 0, 4095, 0, 0),
		(drawing, 1909, 0, 4095, 0, 0),
		(drawing, 1910, 0, 4095, 0, 0),
		(drawing, 1911, 0, 4095, 0, 0),
		(drawing, 1912, 0, 4095, 0, 0),
		(drawing, 1913, 0, 4095, 0, 0),
		(drawing, 1914, 0, 4095, 0, 0),
		(drawing, 1915, 0, 4095, 0, 0),
		(drawing, 1916, 0, 4095, 0, 0),
		(drawing, 1917, 0, 4095, 0, 0),
		(drawing, 1918, 0, 4095, 0, 0),
		(drawing, 1919, 0, 4095, 0, 0),
		(drawing, 1920, 0, 4095, 0, 0),
		(drawing, 1921, 0, 4095, 0, 0),
		(drawing, 1922, 0, 4095, 0, 0),
		(drawing, 1923, 0, 4095, 0, 0),
		(drawing, 1924, 0, 4095, 0, 0),
		(drawing, 1925, 0, 4095, 0, 0),
		(drawing, 1926, 0, 4095, 0, 0),
		(drawing, 1927, 0, 4095, 0, 0),
		(drawing, 1928, 0, 4095, 0, 0),
		(drawing, 1929, 0, 4095, 0, 0),
		(drawing, 1930, 0, 4095, 0, 0),
		(drawing, 1931, 0, 4095, 0, 0),
		(drawing, 1932, 0, 4095, 0, 0),
		(drawing, 1933, 0, 4095, 0, 0),
		(drawing, 1934, 0, 4095, 0, 0),
		(drawing, 1935, 0, 4095, 0, 0),
		(drawing, 1936, 0, 4095, 0, 0),
		(drawing, 1937, 0, 4095, 0, 0),
		(drawing, 1938, 0, 4095, 0, 0),
		(drawing, 1939, 0, 4095, 0, 0),
		(drawing, 1940, 0, 4095, 0, 0),
		(drawing, 1941, 0, 4095, 0, 0),
		(drawing, 1942, 0, 4095, 0, 0),
		(drawing, 1943, 0, 4095, 0, 0),
		(drawing, 1944, 0, 4095, 0, 0),
		(drawing, 1945, 0, 4095, 0, 0),
		(drawing, 1946, 0, 4095, 0, 0),
		(drawing, 1947, 0, 4095, 0, 0),
		(drawing, 1948, 0, 4095, 0, 0),
		(drawing, 1949, 0, 4095, 0, 0),
		(drawing, 1950, 0, 4095, 0, 0),
		(drawing, 1951, 0, 4095, 0, 0),
		(drawing, 1952, 0, 4095, 0, 0),
		(drawing, 1953, 0, 4095, 0, 0),
		(drawing, 1954, 0, 4095, 0, 0),
		(drawing, 1955, 0, 4095, 0, 0),
		(drawing, 1956, 0, 4095, 0, 0),
		(drawing, 1957, 0, 4095, 0, 0),
		(drawing, 1958, 0, 4095, 0, 0),
		(drawing, 1959, 0, 4095, 0, 0),
		(drawing, 1960, 0, 4095, 0, 0),
		(drawing, 1961, 0, 4095, 0, 0),
		(drawing, 1962, 0, 4095, 0, 0),
		(drawing, 1963, 0, 4095, 0, 0),
		(drawing, 1964, 0, 4095, 0, 0),
		(drawing, 1965, 0, 4095, 0, 0),
		(drawing, 1966, 0, 4095, 0, 0),
		(drawing, 1967, 0, 4095, 0, 0),
		(drawing, 1968, 0, 4095, 0, 0),
		(drawing, 1969, 0, 4095, 0, 0),
		(drawing, 1970, 0, 4095, 0, 0),
		(drawing, 1971, 0, 4095, 0, 0),
		(drawing, 1972, 0, 4095, 0, 0),
		(drawing, 1973, 0, 4095, 0, 0),
		(drawing, 1974, 0, 4095, 0, 0),
		(drawing, 1975, 0, 4095, 0, 0),
		(drawing, 1976, 0, 4095, 0, 0),
		(drawing, 1977, 0, 4095, 0, 0),
		(drawing, 1978, 0, 4095, 0, 0),
		(drawing, 1979, 0, 4095, 0, 0),
		(drawing, 1980, 0, 4095, 0, 0),
		(drawing, 1981, 0, 4095, 0, 0),
		(drawing, 1982, 0, 4095, 0, 0),
		(drawing, 1983, 0, 4095, 0, 0),
		(drawing, 1984, 0, 4095, 0, 0),
		(drawing, 1985, 0, 4095, 0, 0),
		(drawing, 1986, 0, 4095, 0, 0),
		(drawing, 1987, 0, 4095, 0, 0),
		(drawing, 1988, 0, 4095, 0, 0),
		(drawing, 1989, 0, 4095, 0, 0),
		(drawing, 1990, 0, 4095, 0, 0),
		(drawing, 1991, 0, 4095, 0, 0),
		(drawing, 1992, 0, 4095, 0, 0),
		(drawing, 1993, 0, 4095, 0, 0),
		(drawing, 1994, 0, 4095, 0, 0),
		(drawing, 1995, 0, 4095, 0, 0),
		(drawing, 1996, 0, 4095, 0, 0),
		(drawing, 1997, 0, 4095, 0, 0),
		(drawing, 1998, 0, 4095, 0, 0),
		(drawing, 1999, 0, 4095, 0, 0),
		(drawing, 2000, 0, 4095, 0, 0),
		(drawing, 2001, 0, 4095, 0, 0),
		(drawing, 2002, 0, 4095, 0, 0),
		(drawing, 2003, 0, 4095, 0, 0),
		(drawing, 2004, 0, 4095, 0, 0),
		(drawing, 2005, 0, 4095, 0, 0),
		(drawing, 2006, 0, 4095, 0, 0),
		(drawing, 2007, 0, 4095, 0, 0),
		(drawing, 2008, 0, 4095, 0, 0),
		(drawing, 2009, 0, 4095, 0, 0),
		(drawing, 2010, 0, 4095, 0, 0),
		(drawing, 2011, 0, 4095, 0, 0),
		(drawing, 2012, 0, 4095, 0, 0),
		(drawing, 2013, 0, 4095, 0, 0),
		(drawing, 2014, 0, 4095, 0, 0),
		(drawing, 2015, 0, 4095, 0, 0),
		(drawing, 2016, 0, 4095, 0, 0),
		(drawing, 2017, 0, 4095, 0, 0),
		(drawing, 2018, 0, 4095, 0, 0),
		(drawing, 2019, 0, 4095, 0, 0),
		(drawing, 2020, 0, 4095, 0, 0),
		(drawing, 2021, 0, 4095, 0, 0),
		(drawing, 2022, 0, 4095, 0, 0),
		(drawing, 2023, 0, 4095, 0, 0),
		(drawing, 2024, 0, 4095, 0, 0),
		(drawing, 2025, 0, 4095, 0, 0),
		(drawing, 2026, 0, 4095, 0, 0),
		(drawing, 2027, 0, 4095, 0, 0),
		(drawing, 2028, 0, 4095, 0, 0),
		(drawing, 2029, 0, 4095, 0, 0),
		(drawing, 2030, 0, 4095, 0, 0),
		(drawing, 2031, 0, 4095, 0, 0),
		(drawing, 2032, 0, 4095, 0, 0),
		(drawing, 2033, 0, 4095, 0, 0),
		(drawing, 2034, 0, 4095, 0, 0),
		(drawing, 2035, 0, 4095, 0, 0),
		(drawing, 2036, 0, 4095, 0, 0),
		(drawing, 2037, 0, 4095, 0, 0),
		(drawing, 2038, 0, 4095, 0, 0),
		(drawing, 2039, 0, 4095, 0, 0),
		(drawing, 2040, 0, 4095, 0, 0),
		(drawing, 2041, 0, 4095, 0, 0),
		(drawing, 2042, 0, 4095, 0, 0),
		(drawing, 2043, 0, 4095, 0, 0),
		(drawing, 2044, 0, 4095, 0, 0),
		(drawing, 2045, 0, 4095, 0, 0),
		(drawing, 2046, 0, 4095, 0, 0),
		(drawing, 2047, 0, 4095, 0, 0),
		(drawing, 2048, 0, 4095, 0, 0),
		(drawing, 2049, 0, 4095, 0, 0),
		(drawing, 2050, 0, 4095, 0, 0),
		(drawing, 2051, 0, 4095, 0, 0),
		(drawing, 2052, 0, 4095, 0, 0),
		(drawing, 2053, 0, 4095, 0, 0),
		(drawing, 2054, 0, 4095, 0, 0),
		(drawing, 2055, 0, 4095, 0, 0),
		(drawing, 2056, 0, 4095, 0, 0),
		(drawing, 2057, 0, 4095, 0, 0),
		(drawing, 2058, 0, 4095, 0, 0),
		(drawing, 2059, 0, 4095, 0, 0),
		(drawing, 2060, 0, 4095, 0, 0),
		(drawing, 2061, 0, 4095, 0, 0),
		(drawing, 2062, 0, 4095, 0, 0),
		(drawing, 2063, 0, 4095, 0, 0),
		(drawing, 2064, 0, 4095, 0, 0),
		(drawing, 2065, 0, 4095, 0, 0),
		(drawing, 2066, 0, 4095, 0, 0),
		(drawing, 2067, 0, 4095, 0, 0),
		(drawing, 2068, 0, 4095, 0, 0),
		(drawing, 2069, 0, 4095, 0, 0),
		(drawing, 2070, 0, 4095, 0, 0),
		(drawing, 2071, 0, 4095, 0, 0),
		(drawing, 2072, 0, 4095, 0, 0),
		(drawing, 2073, 0, 4095, 0, 0),
		(drawing, 2074, 0, 4095, 0, 0),
		(drawing, 2075, 0, 4095, 0, 0),
		(drawing, 2076, 0, 4095, 0, 0),
		(drawing, 2077, 0, 4095, 0, 0),
		(drawing, 2078, 0, 4095, 0, 0),
		(drawing, 2079, 0, 4095, 0, 0),
		(drawing, 2080, 0, 4095, 0, 0),
		(drawing, 2081, 0, 4095, 0, 0),
		(drawing, 2082, 0, 4095, 0, 0),
		(drawing, 2083, 0, 4095, 0, 0),
		(drawing, 2084, 0, 4095, 0, 0),
		(drawing, 2085, 0, 4095, 0, 0),
		(drawing, 2086, 0, 4095, 0, 0),
		(drawing, 2087, 0, 4095, 0, 0),
		(drawing, 2088, 0, 4095, 0, 0),
		(drawing, 2089, 0, 4095, 0, 0),
		(drawing, 2090, 0, 4095, 0, 0),
		(drawing, 2091, 0, 4095, 0, 0),
		(drawing, 2092, 0, 4095, 0, 0),
		(drawing, 2093, 0, 4095, 0, 0),
		(drawing, 2094, 0, 4095, 0, 0),
		(drawing, 2095, 0, 4095, 0, 0),
		(drawing, 2096, 0, 4095, 0, 0),
		(drawing, 2097, 0, 4095, 0, 0),
		(drawing, 2098, 0, 4095, 0, 0),
		(drawing, 2099, 0, 4095, 0, 0),
		(drawing, 2100, 0, 4095, 0, 0),
		(drawing, 2101, 0, 4095, 0, 0),
		(drawing, 2102, 0, 4095, 0, 0),
		(drawing, 2103, 0, 4095, 0, 0),
		(drawing, 2104, 0, 4095, 0, 0),
		(drawing, 2105, 0, 4095, 0, 0),
		(drawing, 2106, 0, 4095, 0, 0),
		(drawing, 2107, 0, 4095, 0, 0),
		(drawing, 2108, 0, 4095, 0, 0),
		(drawing, 2109, 0, 4095, 0, 0),
		(drawing, 2110, 0, 4095, 0, 0),
		(drawing, 2111, 0, 4095, 0, 0),
		(drawing, 2112, 0, 4095, 0, 0),
		(drawing, 2113, 0, 4095, 0, 0),
		(drawing, 2114, 0, 4095, 0, 0),
		(drawing, 2115, 0, 4095, 0, 0),
		(drawing, 2116, 0, 4095, 0, 0),
		(drawing, 2117, 0, 4095, 0, 0),
		(drawing, 2118, 0, 4095, 0, 0),
		(drawing, 2119, 0, 4095, 0, 0),
		(drawing, 2120, 0, 4095, 0, 0),
		(drawing, 2121, 0, 4095, 0, 0),
		(drawing, 2122, 0, 4095, 0, 0),
		(drawing, 2123, 0, 4095, 0, 0),
		(drawing, 2124, 0, 4095, 0, 0),
		(drawing, 2125, 0, 4095, 0, 0),
		(drawing, 2126, 0, 4095, 0, 0),
		(drawing, 2127, 0, 4095, 0, 0),
		(drawing, 2128, 0, 4095, 0, 0),
		(drawing, 2129, 0, 4095, 0, 0),
		(drawing, 2130, 0, 4095, 0, 0),
		(drawing, 2131, 0, 4095, 0, 0),
		(drawing, 2132, 0, 4095, 0, 0),
		(drawing, 2133, 0, 4095, 0, 0),
		(drawing, 2134, 0, 4095, 0, 0),
		(drawing, 2135, 0, 4095, 0, 0),
		(drawing, 2136, 0, 4095, 0, 0),
		(drawing, 2137, 0, 4095, 0, 0),
		(drawing, 2138, 0, 4095, 0, 0),
		(drawing, 2139, 0, 4095, 0, 0),
		(drawing, 2140, 0, 4095, 0, 0),
		(drawing, 2141, 0, 4095, 0, 0),
		(drawing, 2142, 0, 4095, 0, 0),
		(drawing, 2143, 0, 4095, 0, 0),
		(drawing, 2144, 0, 4095, 0, 0),
		(drawing, 2145, 0, 4095, 0, 0),
		(drawing, 2146, 0, 4095, 0, 0),
		(drawing, 2147, 0, 4095, 0, 0),
		(drawing, 2148, 0, 4095, 0, 0),
		(drawing, 2149, 0, 4095, 0, 0),
		(drawing, 2150, 0, 4095, 0, 0),
		(drawing, 2151, 0, 4095, 0, 0),
		(drawing, 2152, 0, 4095, 0, 0),
		(drawing, 2153, 0, 4095, 0, 0),
		(drawing, 2154, 0, 4095, 0, 0),
		(drawing, 2155, 0, 4095, 0, 0),
		(drawing, 2156, 0, 4095, 0, 0),
		(drawing, 2157, 0, 4095, 0, 0),
		(drawing, 2158, 0, 4095, 0, 0),
		(drawing, 2159, 0, 4095, 0, 0),
		(drawing, 2160, 0, 4095, 0, 0),
		(drawing, 2161, 0, 4095, 0, 0),
		(drawing, 2162, 0, 4095, 0, 0),
		(drawing, 2163, 0, 4095, 0, 0),
		(drawing, 2164, 0, 4095, 0, 0),
		(drawing, 2165, 0, 4095, 0, 0),
		(drawing, 2166, 0, 4095, 0, 0),
		(drawing, 2167, 0, 4095, 0, 0),
		(drawing, 2168, 0, 4095, 0, 0),
		(drawing, 2169, 0, 4095, 0, 0),
		(drawing, 2170, 0, 4095, 0, 0),
		(drawing, 2171, 0, 4095, 0, 0),
		(drawing, 2172, 0, 4095, 0, 0),
		(drawing, 2173, 0, 4095, 0, 0),
		(drawing, 2174, 0, 4095, 0, 0),
		(drawing, 2175, 0, 4095, 0, 0),
		(drawing, 2176, 0, 4095, 0, 0),
		(drawing, 2177, 0, 4095, 0, 0),
		(drawing, 2178, 0, 4095, 0, 0),
		(drawing, 2179, 0, 4095, 0, 0),
		(drawing, 2180, 0, 4095, 0, 0),
		(drawing, 2181, 0, 4095, 0, 0),
		(drawing, 2182, 0, 4095, 0, 0),
		(drawing, 2183, 0, 4095, 0, 0),
		(drawing, 2184, 0, 4095, 0, 0),
		(drawing, 2185, 0, 4095, 0, 0),
		(drawing, 2186, 0, 4095, 0, 0),
		(drawing, 2187, 0, 4095, 0, 0),
		(drawing, 2188, 0, 4095, 0, 0),
		(drawing, 2189, 0, 4095, 0, 0),
		(drawing, 2190, 0, 4095, 0, 0),
		(drawing, 2191, 0, 4095, 0, 0),
		(drawing, 2192, 0, 4095, 0, 0),
		(drawing, 2193, 0, 4095, 0, 0),
		(drawing, 2194, 0, 4095, 0, 0),
		(drawing, 2195, 0, 4095, 0, 0),
		(drawing, 2196, 0, 4095, 0, 0),
		(drawing, 2197, 0, 4095, 0, 0),
		(drawing, 2198, 0, 4095, 0, 0),
		(drawing, 2199, 0, 4095, 0, 0),
		(drawing, 2200, 0, 4095, 0, 0),
		(drawing, 2201, 0, 4095, 0, 0),
		(drawing, 2202, 0, 4095, 0, 0),
		(drawing, 2203, 0, 4095, 0, 0),
		(drawing, 2204, 0, 4095, 0, 0),
		(drawing, 2205, 0, 4095, 0, 0),
		(drawing, 2206, 0, 4095, 0, 0),
		(drawing, 2207, 0, 4095, 0, 0),
		(drawing, 2208, 0, 4095, 0, 0),
		(drawing, 2209, 0, 4095, 0, 0),
		(drawing, 2210, 0, 4095, 0, 0),
		(drawing, 2211, 0, 4095, 0, 0),
		(drawing, 2212, 0, 4095, 0, 0),
		(drawing, 2213, 0, 4095, 0, 0),
		(drawing, 2214, 0, 4095, 0, 0),
		(drawing, 2215, 0, 4095, 0, 0),
		(drawing, 2216, 0, 4095, 0, 0),
		(drawing, 2217, 0, 4095, 0, 0),
		(drawing, 2218, 0, 4095, 0, 0),
		(drawing, 2219, 0, 4095, 0, 0),
		(drawing, 2220, 0, 4095, 0, 0),
		(drawing, 2221, 0, 4095, 0, 0),
		(drawing, 2222, 0, 4095, 0, 0),
		(drawing, 2223, 0, 4095, 0, 0),
		(drawing, 2224, 0, 4095, 0, 0),
		(drawing, 2225, 0, 4095, 0, 0),
		(drawing, 2226, 0, 4095, 0, 0),
		(drawing, 2227, 0, 4095, 0, 0),
		(drawing, 2228, 0, 4095, 0, 0),
		(drawing, 2229, 0, 4095, 0, 0),
		(drawing, 2230, 0, 4095, 0, 0),
		(drawing, 2231, 0, 4095, 0, 0),
		(drawing, 2232, 0, 4095, 0, 0),
		(drawing, 2233, 0, 4095, 0, 0),
		(drawing, 2234, 0, 4095, 0, 0),
		(drawing, 2235, 0, 4095, 0, 0),
		(drawing, 2236, 0, 4095, 0, 0),
		(drawing, 2237, 0, 4095, 0, 0),
		(drawing, 2238, 0, 4095, 0, 0),
		(drawing, 2239, 0, 4095, 0, 0),
		(drawing, 2240, 0, 4095, 0, 0),
		(drawing, 2241, 0, 4095, 0, 0),
		(drawing, 2242, 0, 4095, 0, 0),
		(drawing, 2243, 0, 4095, 0, 0),
		(drawing, 2244, 0, 4095, 0, 0),
		(drawing, 2245, 0, 4095, 0, 0),
		(drawing, 2246, 0, 4095, 0, 0),
		(drawing, 2247, 0, 4095, 0, 0),
		(drawing, 2248, 0, 4095, 0, 0),
		(drawing, 2249, 0, 4095, 0, 0),
		(drawing, 2250, 0, 4095, 0, 0),
		(drawing, 2251, 0, 4095, 0, 0),
		(drawing, 2252, 0, 4095, 0, 0),
		(drawing, 2253, 0, 4095, 0, 0),
		(drawing, 2254, 0, 4095, 0, 0),
		(drawing, 2255, 0, 4095, 0, 0),
		(drawing, 2256, 0, 4095, 0, 0),
		(drawing, 2257, 0, 4095, 0, 0),
		(drawing, 2258, 0, 4095, 0, 0),
		(drawing, 2259, 0, 4095, 0, 0),
		(drawing, 2260, 0, 4095, 0, 0),
		(drawing, 2261, 0, 4095, 0, 0),
		(drawing, 2262, 0, 4095, 0, 0),
		(drawing, 2263, 0, 4095, 0, 0),
		(drawing, 2264, 0, 4095, 0, 0),
		(drawing, 2265, 0, 4095, 0, 0),
		(drawing, 2266, 0, 4095, 0, 0),
		(drawing, 2267, 0, 4095, 0, 0),
		(drawing, 2268, 0, 4095, 0, 0),
		(drawing, 2269, 0, 4095, 0, 0),
		(drawing, 2270, 0, 4095, 0, 0),
		(drawing, 2271, 0, 4095, 0, 0),
		(drawing, 2272, 0, 4095, 0, 0),
		(drawing, 2273, 0, 4095, 0, 0),
		(drawing, 2274, 0, 4095, 0, 0),
		(drawing, 2275, 0, 4095, 0, 0),
		(drawing, 2276, 0, 4095, 0, 0),
		(drawing, 2277, 0, 4095, 0, 0),
		(drawing, 2278, 0, 4095, 0, 0),
		(drawing, 2279, 0, 4095, 0, 0),
		(drawing, 2280, 0, 4095, 0, 0),
		(drawing, 2281, 0, 4095, 0, 0),
		(drawing, 2282, 0, 4095, 0, 0),
		(drawing, 2283, 0, 4095, 0, 0),
		(drawing, 2284, 0, 4095, 0, 0),
		(drawing, 2285, 0, 4095, 0, 0),
		(drawing, 2286, 0, 4095, 0, 0),
		(drawing, 2287, 0, 4095, 0, 0),
		(drawing, 2288, 0, 4095, 0, 0),
		(drawing, 2289, 0, 4095, 0, 0),
		(drawing, 2290, 0, 4095, 0, 0),
		(drawing, 2291, 0, 4095, 0, 0),
		(drawing, 2292, 0, 4095, 0, 0),
		(drawing, 2293, 0, 4095, 0, 0),
		(drawing, 2294, 0, 4095, 0, 0),
		(drawing, 2295, 0, 4095, 0, 0),
		(drawing, 2296, 0, 4095, 0, 0),
		(drawing, 2297, 0, 4095, 0, 0),
		(drawing, 2298, 0, 4095, 0, 0),
		(drawing, 2299, 0, 4095, 0, 0),
		(drawing, 2300, 0, 4095, 0, 0),
		(drawing, 2301, 0, 4095, 0, 0),
		(drawing, 2302, 0, 4095, 0, 0),
		(drawing, 2303, 0, 4095, 0, 0),
		(drawing, 2304, 0, 4095, 0, 0),
		(drawing, 2305, 0, 4095, 0, 0),
		(drawing, 2306, 0, 4095, 0, 0),
		(drawing, 2307, 0, 4095, 0, 0),
		(drawing, 2308, 0, 4095, 0, 0),
		(drawing, 2309, 0, 4095, 0, 0),
		(drawing, 2310, 0, 4095, 0, 0),
		(drawing, 2311, 0, 4095, 0, 0),
		(drawing, 2312, 0, 4095, 0, 0),
		(drawing, 2313, 0, 4095, 0, 0),
		(drawing, 2314, 0, 4095, 0, 0),
		(drawing, 2315, 0, 4095, 0, 0),
		(drawing, 2316, 0, 4095, 0, 0),
		(drawing, 2317, 0, 4095, 0, 0),
		(drawing, 2318, 0, 4095, 0, 0),
		(drawing, 2319, 0, 4095, 0, 0),
		(drawing, 2320, 0, 4095, 0, 0),
		(drawing, 2321, 0, 4095, 0, 0),
		(drawing, 2322, 0, 4095, 0, 0),
		(drawing, 2323, 0, 4095, 0, 0),
		(drawing, 2324, 0, 4095, 0, 0),
		(drawing, 2325, 0, 4095, 0, 0),
		(drawing, 2326, 0, 4095, 0, 0),
		(drawing, 2327, 0, 4095, 0, 0),
		(drawing, 2328, 0, 4095, 0, 0),
		(drawing, 2329, 0, 4095, 0, 0),
		(drawing, 2330, 0, 4095, 0, 0),
		(drawing, 2331, 0, 4095, 0, 0),
		(drawing, 2332, 0, 4095, 0, 0),
		(drawing, 2333, 0, 4095, 0, 0),
		(drawing, 2334, 0, 4095, 0, 0),
		(drawing, 2335, 0, 4095, 0, 0),
		(drawing, 2336, 0, 4095, 0, 0),
		(drawing, 2337, 0, 4095, 0, 0),
		(drawing, 2338, 0, 4095, 0, 0),
		(drawing, 2339, 0, 4095, 0, 0),
		(drawing, 2340, 0, 4095, 0, 0),
		(drawing, 2341, 0, 4095, 0, 0),
		(drawing, 2342, 0, 4095, 0, 0),
		(drawing, 2343, 0, 4095, 0, 0),
		(drawing, 2344, 0, 4095, 0, 0),
		(drawing, 2345, 0, 4095, 0, 0),
		(drawing, 2346, 0, 4095, 0, 0),
		(drawing, 2347, 0, 4095, 0, 0),
		(drawing, 2348, 0, 4095, 0, 0),
		(drawing, 2349, 0, 4095, 0, 0),
		(drawing, 2350, 0, 4095, 0, 0),
		(drawing, 2351, 0, 4095, 0, 0),
		(drawing, 2352, 0, 4095, 0, 0),
		(drawing, 2353, 0, 4095, 0, 0),
		(drawing, 2354, 0, 4095, 0, 0),
		(drawing, 2355, 0, 4095, 0, 0),
		(drawing, 2356, 0, 4095, 0, 0),
		(drawing, 2357, 0, 4095, 0, 0),
		(drawing, 2358, 0, 4095, 0, 0),
		(drawing, 2359, 0, 4095, 0, 0),
		(drawing, 2360, 0, 4095, 0, 0),
		(drawing, 2361, 0, 4095, 0, 0),
		(drawing, 2362, 0, 4095, 0, 0),
		(drawing, 2363, 0, 4095, 0, 0),
		(drawing, 2364, 0, 4095, 0, 0),
		(drawing, 2365, 0, 4095, 0, 0),
		(drawing, 2366, 0, 4095, 0, 0),
		(drawing, 2367, 0, 4095, 0, 0),
		(drawing, 2368, 0, 4095, 0, 0),
		(drawing, 2369, 0, 4095, 0, 0),
		(drawing, 2370, 0, 4095, 0, 0),
		(drawing, 2371, 0, 4095, 0, 0),
		(drawing, 2372, 0, 4095, 0, 0),
		(drawing, 2373, 0, 4095, 0, 0),
		(drawing, 2374, 0, 4095, 0, 0),
		(drawing, 2375, 0, 4095, 0, 0),
		(drawing, 2376, 0, 4095, 0, 0),
		(drawing, 2377, 0, 4095, 0, 0),
		(drawing, 2378, 0, 4095, 0, 0),
		(drawing, 2379, 0, 4095, 0, 0),
		(drawing, 2380, 0, 4095, 0, 0),
		(drawing, 2381, 0, 4095, 0, 0),
		(drawing, 2382, 0, 4095, 0, 0),
		(drawing, 2383, 0, 4095, 0, 0),
		(drawing, 2384, 0, 4095, 0, 0),
		(drawing, 2385, 0, 4095, 0, 0),
		(drawing, 2386, 0, 4095, 0, 0),
		(drawing, 2387, 0, 4095, 0, 0),
		(drawing, 2388, 0, 4095, 0, 0),
		(drawing, 2389, 0, 4095, 0, 0),
		(drawing, 2390, 0, 4095, 0, 0),
		(drawing, 2391, 0, 4095, 0, 0),
		(drawing, 2392, 0, 4095, 0, 0),
		(drawing, 2393, 0, 4095, 0, 0),
		(drawing, 2394, 0, 4095, 0, 0),
		(drawing, 2395, 0, 4095, 0, 0),
		(drawing, 2396, 0, 4095, 0, 0),
		(drawing, 2397, 0, 4095, 0, 0),
		(drawing, 2398, 0, 4095, 0, 0),
		(drawing, 2399, 0, 4095, 0, 0),
		(drawing, 2400, 0, 4095, 0, 0),
		(drawing, 2401, 0, 4095, 0, 0),
		(drawing, 2402, 0, 4095, 0, 0),
		(drawing, 2403, 0, 4095, 0, 0),
		(drawing, 2404, 0, 4095, 0, 0),
		(drawing, 2405, 0, 4095, 0, 0),
		(drawing, 2406, 0, 4095, 0, 0),
		(drawing, 2407, 0, 4095, 0, 0),
		(drawing, 2408, 0, 4095, 0, 0),
		(drawing, 2409, 0, 4095, 0, 0),
		(drawing, 2410, 0, 4095, 0, 0),
		(drawing, 2411, 0, 4095, 0, 0),
		(drawing, 2412, 0, 4095, 0, 0),
		(drawing, 2413, 0, 4095, 0, 0),
		(drawing, 2414, 0, 4095, 0, 0),
		(drawing, 2415, 0, 4095, 0, 0),
		(drawing, 2416, 0, 4095, 0, 0),
		(drawing, 2417, 0, 4095, 0, 0),
		(drawing, 2418, 0, 4095, 0, 0),
		(drawing, 2419, 0, 4095, 0, 0),
		(drawing, 2420, 0, 4095, 0, 0),
		(drawing, 2421, 0, 4095, 0, 0),
		(drawing, 2422, 0, 4095, 0, 0),
		(drawing, 2423, 0, 4095, 0, 0),
		(drawing, 2424, 0, 4095, 0, 0),
		(drawing, 2425, 0, 4095, 0, 0),
		(drawing, 2426, 0, 4095, 0, 0),
		(drawing, 2427, 0, 4095, 0, 0),
		(drawing, 2428, 0, 4095, 0, 0),
		(drawing, 2429, 0, 4095, 0, 0),
		(drawing, 2430, 0, 4095, 0, 0),
		(drawing, 2431, 0, 4095, 0, 0),
		(drawing, 2432, 0, 4095, 0, 0),
		(drawing, 2433, 0, 4095, 0, 0),
		(drawing, 2434, 0, 4095, 0, 0),
		(drawing, 2435, 0, 4095, 0, 0),
		(drawing, 2436, 0, 4095, 0, 0),
		(drawing, 2437, 0, 4095, 0, 0),
		(drawing, 2438, 0, 4095, 0, 0),
		(drawing, 2439, 0, 4095, 0, 0),
		(drawing, 2440, 0, 4095, 0, 0),
		(drawing, 2441, 0, 4095, 0, 0),
		(drawing, 2442, 0, 4095, 0, 0),
		(drawing, 2443, 0, 4095, 0, 0),
		(drawing, 2444, 0, 4095, 0, 0),
		(drawing, 2445, 0, 4095, 0, 0),
		(drawing, 2446, 0, 4095, 0, 0),
		(drawing, 2447, 0, 4095, 0, 0),
		(drawing, 2448, 0, 4095, 0, 0),
		(drawing, 2449, 0, 4095, 0, 0),
		(drawing, 2450, 0, 4095, 0, 0),
		(drawing, 2451, 0, 4095, 0, 0),
		(drawing, 2452, 0, 4095, 0, 0),
		(drawing, 2453, 0, 4095, 0, 0),
		(drawing, 2454, 0, 4095, 0, 0),
		(drawing, 2455, 0, 4095, 0, 0),
		(drawing, 2456, 0, 4095, 0, 0),
		(drawing, 2457, 0, 4095, 0, 0),
		(drawing, 2458, 0, 4095, 0, 0),
		(drawing, 2459, 0, 4095, 0, 0),
		(drawing, 2460, 0, 4095, 0, 0),
		(drawing, 2461, 0, 4095, 0, 0),
		(drawing, 2462, 0, 4095, 0, 0),
		(drawing, 2463, 0, 4095, 0, 0),
		(drawing, 2464, 0, 4095, 0, 0),
		(drawing, 2465, 0, 4095, 0, 0),
		(drawing, 2466, 0, 4095, 0, 0),
		(drawing, 2467, 0, 4095, 0, 0),
		(drawing, 2468, 0, 4095, 0, 0),
		(drawing, 2469, 0, 4095, 0, 0),
		(drawing, 2470, 0, 4095, 0, 0),
		(drawing, 2471, 0, 4095, 0, 0),
		(drawing, 2472, 0, 4095, 0, 0),
		(drawing, 2473, 0, 4095, 0, 0),
		(drawing, 2474, 0, 4095, 0, 0),
		(drawing, 2475, 0, 4095, 0, 0),
		(drawing, 2476, 0, 4095, 0, 0),
		(drawing, 2477, 0, 4095, 0, 0),
		(drawing, 2478, 0, 4095, 0, 0),
		(drawing, 2479, 0, 4095, 0, 0),
		(drawing, 2480, 0, 4095, 0, 0),
		(drawing, 2481, 0, 4095, 0, 0),
		(drawing, 2482, 0, 4095, 0, 0),
		(drawing, 2483, 0, 4095, 0, 0),
		(drawing, 2484, 0, 4095, 0, 0),
		(drawing, 2485, 0, 4095, 0, 0),
		(drawing, 2486, 0, 4095, 0, 0),
		(drawing, 2487, 0, 4095, 0, 0),
		(drawing, 2488, 0, 4095, 0, 0),
		(drawing, 2489, 0, 4095, 0, 0),
		(drawing, 2490, 0, 4095, 0, 0),
		(drawing, 2491, 0, 4095, 0, 0),
		(drawing, 2492, 0, 4095, 0, 0),
		(drawing, 2493, 0, 4095, 0, 0),
		(drawing, 2494, 0, 4095, 0, 0),
		(drawing, 2495, 0, 4095, 0, 0),
		(drawing, 2496, 0, 4095, 0, 0),
		(drawing, 2497, 0, 4095, 0, 0),
		(drawing, 2498, 0, 4095, 0, 0),
		(drawing, 2499, 0, 4095, 0, 0),
		(drawing, 2500, 0, 4095, 0, 0),
		(drawing, 2501, 0, 4095, 0, 0),
		(drawing, 2502, 0, 4095, 0, 0),
		(drawing, 2503, 0, 4095, 0, 0),
		(drawing, 2504, 0, 4095, 0, 0),
		(drawing, 2505, 0, 4095, 0, 0),
		(drawing, 2506, 0, 4095, 0, 0),
		(drawing, 2507, 0, 4095, 0, 0),
		(drawing, 2508, 0, 4095, 0, 0),
		(drawing, 2509, 0, 4095, 0, 0),
		(drawing, 2510, 0, 4095, 0, 0),
		(drawing, 2511, 0, 4095, 0, 0),
		(drawing, 2512, 0, 4095, 0, 0),
		(drawing, 2513, 0, 4095, 0, 0),
		(drawing, 2514, 0, 4095, 0, 0),
		(drawing, 2515, 0, 4095, 0, 0),
		(drawing, 2516, 0, 4095, 0, 0),
		(drawing, 2517, 0, 4095, 0, 0),
		(drawing, 2518, 0, 4095, 0, 0),
		(drawing, 2519, 0, 4095, 0, 0),
		(drawing, 2520, 0, 4095, 0, 0),
		(drawing, 2521, 0, 4095, 0, 0),
		(drawing, 2522, 0, 4095, 0, 0),
		(drawing, 2523, 0, 4095, 0, 0),
		(drawing, 2524, 0, 4095, 0, 0),
		(drawing, 2525, 0, 4095, 0, 0),
		(drawing, 2526, 0, 4095, 0, 0),
		(drawing, 2527, 0, 4095, 0, 0),
		(drawing, 2528, 0, 4095, 0, 0),
		(drawing, 2529, 0, 4095, 0, 0),
		(drawing, 2530, 0, 4095, 0, 0),
		(drawing, 2531, 0, 4095, 0, 0),
		(drawing, 2532, 0, 4095, 0, 0),
		(drawing, 2533, 0, 4095, 0, 0),
		(drawing, 2534, 0, 4095, 0, 0),
		(drawing, 2535, 0, 4095, 0, 0),
		(drawing, 2536, 0, 4095, 0, 0),
		(drawing, 2537, 0, 4095, 0, 0),
		(drawing, 2538, 0, 4095, 0, 0),
		(drawing, 2539, 0, 4095, 0, 0),
		(drawing, 2540, 0, 4095, 0, 0),
		(drawing, 2541, 0, 4095, 0, 0),
		(drawing, 2542, 0, 4095, 0, 0),
		(drawing, 2543, 0, 4095, 0, 0),
		(drawing, 2544, 0, 4095, 0, 0),
		(drawing, 2545, 0, 4095, 0, 0),
		(drawing, 2546, 0, 4095, 0, 0),
		(drawing, 2547, 0, 4095, 0, 0),
		(drawing, 2548, 0, 4095, 0, 0),
		(drawing, 2549, 0, 4095, 0, 0),
		(drawing, 2550, 0, 4095, 0, 0),
		(drawing, 2551, 0, 4095, 0, 0),
		(drawing, 2552, 0, 4095, 0, 0),
		(drawing, 2553, 0, 4095, 0, 0),
		(drawing, 2554, 0, 4095, 0, 0),
		(drawing, 2555, 0, 4095, 0, 0),
		(drawing, 2556, 0, 4095, 0, 0),
		(drawing, 2557, 0, 4095, 0, 0),
		(drawing, 2558, 0, 4095, 0, 0),
		(drawing, 2559, 0, 4095, 0, 0),
		(drawing, 2560, 0, 4095, 0, 0),
		(drawing, 2561, 0, 4095, 0, 0),
		(drawing, 2562, 0, 4095, 0, 0),
		(drawing, 2563, 0, 4095, 0, 0),
		(drawing, 2564, 0, 4095, 0, 0),
		(drawing, 2565, 0, 4095, 0, 0),
		(drawing, 2566, 0, 4095, 0, 0),
		(drawing, 2567, 0, 4095, 0, 0),
		(drawing, 2568, 0, 4095, 0, 0),
		(drawing, 2569, 0, 4095, 0, 0),
		(drawing, 2570, 0, 4095, 0, 0),
		(drawing, 2571, 0, 4095, 0, 0),
		(drawing, 2572, 0, 4095, 0, 0),
		(drawing, 2573, 0, 4095, 0, 0),
		(drawing, 2574, 0, 4095, 0, 0),
		(drawing, 2575, 0, 4095, 0, 0),
		(drawing, 2576, 0, 4095, 0, 0),
		(drawing, 2577, 0, 4095, 0, 0),
		(drawing, 2578, 0, 4095, 0, 0),
		(drawing, 2579, 0, 4095, 0, 0),
		(drawing, 2580, 0, 4095, 0, 0),
		(drawing, 2581, 0, 4095, 0, 0),
		(drawing, 2582, 0, 4095, 0, 0),
		(drawing, 2583, 0, 4095, 0, 0),
		(drawing, 2584, 0, 4095, 0, 0),
		(drawing, 2585, 0, 4095, 0, 0),
		(drawing, 2586, 0, 4095, 0, 0),
		(drawing, 2587, 0, 4095, 0, 0),
		(drawing, 2588, 0, 4095, 0, 0),
		(drawing, 2589, 0, 4095, 0, 0),
		(drawing, 2590, 0, 4095, 0, 0),
		(drawing, 2591, 0, 4095, 0, 0),
		(drawing, 2592, 0, 4095, 0, 0),
		(drawing, 2593, 0, 4095, 0, 0),
		(drawing, 2594, 0, 4095, 0, 0),
		(drawing, 2595, 0, 4095, 0, 0),
		(drawing, 2596, 0, 4095, 0, 0),
		(drawing, 2597, 0, 4095, 0, 0),
		(drawing, 2598, 0, 4095, 0, 0),
		(drawing, 2599, 0, 4095, 0, 0),
		(drawing, 2600, 0, 4095, 0, 0),
		(drawing, 2601, 0, 4095, 0, 0),
		(drawing, 2602, 0, 4095, 0, 0),
		(drawing, 2603, 0, 4095, 0, 0),
		(drawing, 2604, 0, 4095, 0, 0),
		(drawing, 2605, 0, 4095, 0, 0),
		(drawing, 2606, 0, 4095, 0, 0),
		(drawing, 2607, 0, 4095, 0, 0),
		(drawing, 2608, 0, 4095, 0, 0),
		(drawing, 2609, 0, 4095, 0, 0),
		(drawing, 2610, 0, 4095, 0, 0),
		(drawing, 2611, 0, 4095, 0, 0),
		(drawing, 2612, 0, 4095, 0, 0),
		(drawing, 2613, 0, 4095, 0, 0),
		(drawing, 2614, 0, 4095, 0, 0),
		(drawing, 2615, 0, 4095, 0, 0),
		(drawing, 2616, 0, 4095, 0, 0),
		(drawing, 2617, 0, 4095, 0, 0),
		(drawing, 2618, 0, 4095, 0, 0),
		(drawing, 2619, 0, 4095, 0, 0),
		(drawing, 2620, 0, 4095, 0, 0),
		(drawing, 2621, 0, 4095, 0, 0),
		(drawing, 2622, 0, 4095, 0, 0),
		(drawing, 2623, 0, 4095, 0, 0),
		(drawing, 2624, 0, 4095, 0, 0),
		(drawing, 2625, 0, 4095, 0, 0),
		(drawing, 2626, 0, 4095, 0, 0),
		(drawing, 2627, 0, 4095, 0, 0),
		(drawing, 2628, 0, 4095, 0, 0),
		(drawing, 2629, 0, 4095, 0, 0),
		(drawing, 2630, 0, 4095, 0, 0),
		(drawing, 2631, 0, 4095, 0, 0),
		(drawing, 2632, 0, 4095, 0, 0),
		(drawing, 2633, 0, 4095, 0, 0),
		(drawing, 2634, 0, 4095, 0, 0),
		(drawing, 2635, 0, 4095, 0, 0),
		(drawing, 2636, 0, 4095, 0, 0),
		(drawing, 2637, 0, 4095, 0, 0),
		(drawing, 2638, 0, 4095, 0, 0),
		(drawing, 2639, 0, 4095, 0, 0),
		(drawing, 2640, 0, 4095, 0, 0),
		(drawing, 2641, 0, 4095, 0, 0),
		(drawing, 2642, 0, 4095, 0, 0),
		(drawing, 2643, 0, 4095, 0, 0),
		(drawing, 2644, 0, 4095, 0, 0),
		(drawing, 2645, 0, 4095, 0, 0),
		(drawing, 2646, 0, 4095, 0, 0),
		(drawing, 2647, 0, 4095, 0, 0),
		(drawing, 2648, 0, 4095, 0, 0),
		(drawing, 2649, 0, 4095, 0, 0),
		(drawing, 2650, 0, 4095, 0, 0),
		(drawing, 2651, 0, 4095, 0, 0),
		(drawing, 2652, 0, 4095, 0, 0),
		(drawing, 2653, 0, 4095, 0, 0),
		(drawing, 2654, 0, 4095, 0, 0),
		(drawing, 2655, 0, 4095, 0, 0),
		(drawing, 2656, 0, 4095, 0, 0),
		(drawing, 2657, 0, 4095, 0, 0),
		(drawing, 2658, 0, 4095, 0, 0),
		(drawing, 2659, 0, 4095, 0, 0),
		(drawing, 2660, 0, 4095, 0, 0),
		(drawing, 2661, 0, 4095, 0, 0),
		(drawing, 2662, 0, 4095, 0, 0),
		(drawing, 2663, 0, 4095, 0, 0),
		(drawing, 2664, 0, 4095, 0, 0),
		(drawing, 2665, 0, 4095, 0, 0),
		(drawing, 2666, 0, 4095, 0, 0),
		(drawing, 2667, 0, 4095, 0, 0),
		(drawing, 2668, 0, 4095, 0, 0),
		(drawing, 2669, 0, 4095, 0, 0),
		(drawing, 2670, 0, 4095, 0, 0),
		(drawing, 2671, 0, 4095, 0, 0),
		(drawing, 2672, 0, 4095, 0, 0),
		(drawing, 2673, 0, 4095, 0, 0),
		(drawing, 2674, 0, 4095, 0, 0),
		(drawing, 2675, 0, 4095, 0, 0),
		(drawing, 2676, 0, 4095, 0, 0),
		(drawing, 2677, 0, 4095, 0, 0),
		(drawing, 2678, 0, 4095, 0, 0),
		(drawing, 2679, 0, 4095, 0, 0),
		(drawing, 2680, 0, 4095, 0, 0),
		(drawing, 2681, 0, 4095, 0, 0),
		(drawing, 2682, 0, 4095, 0, 0),
		(drawing, 2683, 0, 4095, 0, 0),
		(drawing, 2684, 0, 4095, 0, 0),
		(drawing, 2685, 0, 4095, 0, 0),
		(drawing, 2686, 0, 4095, 0, 0),
		(drawing, 2687, 0, 4095, 0, 0),
		(drawing, 2688, 0, 4095, 0, 0),
		(drawing, 2689, 0, 4095, 0, 0),
		(drawing, 2690, 0, 4095, 0, 0),
		(drawing, 2691, 0, 4095, 0, 0),
		(drawing, 2692, 0, 4095, 0, 0),
		(drawing, 2693, 0, 4095, 0, 0),
		(drawing, 2694, 0, 4095, 0, 0),
		(drawing, 2695, 0, 4095, 0, 0),
		(drawing, 2696, 0, 4095, 0, 0),
		(drawing, 2697, 0, 4095, 0, 0),
		(drawing, 2698, 0, 4095, 0, 0),
		(drawing, 2699, 0, 4095, 0, 0),
		(drawing, 2700, 0, 4095, 0, 0),
		(drawing, 2701, 0, 4095, 0, 0),
		(drawing, 2702, 0, 4095, 0, 0),
		(drawing, 2703, 0, 4095, 0, 0),
		(drawing, 2704, 0, 4095, 0, 0),
		(drawing, 2705, 0, 4095, 0, 0),
		(drawing, 2706, 0, 4095, 0, 0),
		(drawing, 2707, 0, 4095, 0, 0),
		(drawing, 2708, 0, 4095, 0, 0),
		(drawing, 2709, 0, 4095, 0, 0),
		(drawing, 2710, 0, 4095, 0, 0),
		(drawing, 2711, 0, 4095, 0, 0),
		(drawing, 2712, 0, 4095, 0, 0),
		(drawing, 2713, 0, 4095, 0, 0),
		(drawing, 2714, 0, 4095, 0, 0),
		(drawing, 2715, 0, 4095, 0, 0),
		(drawing, 2716, 0, 4095, 0, 0),
		(drawing, 2717, 0, 4095, 0, 0),
		(drawing, 2718, 0, 4095, 0, 0),
		(drawing, 2719, 0, 4095, 0, 0),
		(drawing, 2720, 0, 4095, 0, 0),
		(drawing, 2721, 0, 4095, 0, 0),
		(drawing, 2722, 0, 4095, 0, 0),
		(drawing, 2723, 0, 4095, 0, 0),
		(drawing, 2724, 0, 4095, 0, 0),
		(drawing, 2725, 0, 4095, 0, 0),
		(drawing, 2726, 0, 4095, 0, 0),
		(drawing, 2727, 0, 4095, 0, 0),
		(drawing, 2728, 0, 4095, 0, 0),
		(drawing, 2729, 0, 4095, 0, 0),
		(drawing, 2730, 0, 4095, 0, 0),
		(drawing, 2731, 0, 4095, 0, 0),
		(drawing, 2732, 0, 4095, 0, 0),
		(drawing, 2733, 0, 4095, 0, 0),
		(drawing, 2734, 0, 4095, 0, 0),
		(drawing, 2735, 0, 4095, 0, 0),
		(drawing, 2736, 0, 4095, 0, 0),
		(drawing, 2737, 0, 4095, 0, 0),
		(drawing, 2738, 0, 4095, 0, 0),
		(drawing, 2739, 0, 4095, 0, 0),
		(drawing, 2740, 0, 4095, 0, 0),
		(drawing, 2741, 0, 4095, 0, 0),
		(drawing, 2742, 0, 4095, 0, 0),
		(drawing, 2743, 0, 4095, 0, 0),
		(drawing, 2744, 0, 4095, 0, 0),
		(drawing, 2745, 0, 4095, 0, 0),
		(drawing, 2746, 0, 4095, 0, 0),
		(drawing, 2747, 0, 4095, 0, 0),
		(drawing, 2748, 0, 4095, 0, 0),
		(drawing, 2749, 0, 4095, 0, 0),
		(drawing, 2750, 0, 4095, 0, 0),
		(drawing, 2751, 0, 4095, 0, 0),
		(drawing, 2752, 0, 4095, 0, 0),
		(drawing, 2753, 0, 4095, 0, 0),
		(drawing, 2754, 0, 4095, 0, 0),
		(drawing, 2755, 0, 4095, 0, 0),
		(drawing, 2756, 0, 4095, 0, 0),
		(drawing, 2757, 0, 4095, 0, 0),
		(drawing, 2758, 0, 4095, 0, 0),
		(drawing, 2759, 0, 4095, 0, 0),
		(drawing, 2760, 0, 4095, 0, 0),
		(drawing, 2761, 0, 4095, 0, 0),
		(drawing, 2762, 0, 4095, 0, 0),
		(drawing, 2763, 0, 4095, 0, 0),
		(drawing, 2764, 0, 4095, 0, 0),
		(drawing, 2765, 0, 4095, 0, 0),
		(drawing, 2766, 0, 4095, 0, 0),
		(drawing, 2767, 0, 4095, 0, 0),
		(drawing, 2768, 0, 4095, 0, 0),
		(drawing, 2769, 0, 4095, 0, 0),
		(drawing, 2770, 0, 4095, 0, 0),
		(drawing, 2771, 0, 4095, 0, 0),
		(drawing, 2772, 0, 4095, 0, 0),
		(drawing, 2773, 0, 4095, 0, 0),
		(drawing, 2774, 0, 4095, 0, 0),
		(drawing, 2775, 0, 4095, 0, 0),
		(drawing, 2776, 0, 4095, 0, 0),
		(drawing, 2777, 0, 4095, 0, 0),
		(drawing, 2778, 0, 4095, 0, 0),
		(drawing, 2779, 0, 4095, 0, 0),
		(drawing, 2780, 0, 4095, 0, 0),
		(drawing, 2781, 0, 4095, 0, 0),
		(drawing, 2782, 0, 4095, 0, 0),
		(drawing, 2783, 0, 4095, 0, 0),
		(drawing, 2784, 0, 4095, 0, 0),
		(drawing, 2785, 0, 4095, 0, 0),
		(drawing, 2786, 0, 4095, 0, 0),
		(drawing, 2787, 0, 4095, 0, 0),
		(drawing, 2788, 0, 4095, 0, 0),
		(drawing, 2789, 0, 4095, 0, 0),
		(drawing, 2790, 0, 4095, 0, 0),
		(drawing, 2791, 0, 4095, 0, 0),
		(drawing, 2792, 0, 4095, 0, 0),
		(drawing, 2793, 0, 4095, 0, 0),
		(drawing, 2794, 0, 4095, 0, 0),
		(drawing, 2795, 0, 4095, 0, 0),
		(drawing, 2796, 0, 4095, 0, 0),
		(drawing, 2797, 0, 4095, 0, 0),
		(drawing, 2798, 0, 4095, 0, 0),
		(drawing, 2799, 0, 4095, 0, 0),
		(drawing, 2800, 0, 4095, 0, 0),
		(drawing, 2801, 0, 4095, 0, 0),
		(drawing, 2802, 0, 4095, 0, 0),
		(drawing, 2803, 0, 4095, 0, 0),
		(drawing, 2804, 0, 4095, 0, 0),
		(drawing, 2805, 0, 4095, 0, 0),
		(drawing, 2806, 0, 4095, 0, 0),
		(drawing, 2807, 0, 4095, 0, 0),
		(drawing, 2808, 0, 4095, 0, 0),
		(drawing, 2809, 0, 4095, 0, 0),
		(drawing, 2810, 0, 4095, 0, 0),
		(drawing, 2811, 0, 4095, 0, 0),
		(drawing, 2812, 0, 4095, 0, 0),
		(drawing, 2813, 0, 4095, 0, 0),
		(drawing, 2814, 0, 4095, 0, 0),
		(drawing, 2815, 0, 4095, 0, 0),
		(drawing, 2816, 0, 4095, 0, 0),
		(drawing, 2817, 0, 4095, 0, 0),
		(drawing, 2818, 0, 4095, 0, 0),
		(drawing, 2819, 0, 4095, 0, 0),
		(drawing, 2820, 0, 4095, 0, 0),
		(drawing, 2821, 0, 4095, 0, 0),
		(drawing, 2822, 0, 4095, 0, 0),
		(drawing, 2823, 0, 4095, 0, 0),
		(drawing, 2824, 0, 4095, 0, 0),
		(drawing, 2825, 0, 4095, 0, 0),
		(drawing, 2826, 0, 4095, 0, 0),
		(drawing, 2827, 0, 4095, 0, 0),
		(drawing, 2828, 0, 4095, 0, 0),
		(drawing, 2829, 0, 4095, 0, 0),
		(drawing, 2830, 0, 4095, 0, 0),
		(drawing, 2831, 0, 4095, 0, 0),
		(drawing, 2832, 0, 4095, 0, 0),
		(drawing, 2833, 0, 4095, 0, 0),
		(drawing, 2834, 0, 4095, 0, 0),
		(drawing, 2835, 0, 4095, 0, 0),
		(drawing, 2836, 0, 4095, 0, 0),
		(drawing, 2837, 0, 4095, 0, 0),
		(drawing, 2838, 0, 4095, 0, 0),
		(drawing, 2839, 0, 4095, 0, 0),
		(drawing, 2840, 0, 4095, 0, 0),
		(drawing, 2841, 0, 4095, 0, 0),
		(drawing, 2842, 0, 4095, 0, 0),
		(drawing, 2843, 0, 4095, 0, 0),
		(drawing, 2844, 0, 4095, 0, 0),
		(drawing, 2845, 0, 4095, 0, 0),
		(drawing, 2846, 0, 4095, 0, 0),
		(drawing, 2847, 0, 4095, 0, 0),
		(drawing, 2848, 0, 4095, 0, 0),
		(drawing, 2849, 0, 4095, 0, 0),
		(drawing, 2850, 0, 4095, 0, 0),
		(drawing, 2851, 0, 4095, 0, 0),
		(drawing, 2852, 0, 4095, 0, 0),
		(drawing, 2853, 0, 4095, 0, 0),
		(drawing, 2854, 0, 4095, 0, 0),
		(drawing, 2855, 0, 4095, 0, 0),
		(drawing, 2856, 0, 4095, 0, 0),
		(drawing, 2857, 0, 4095, 0, 0),
		(drawing, 2858, 0, 4095, 0, 0),
		(drawing, 2859, 0, 4095, 0, 0),
		(drawing, 2860, 0, 4095, 0, 0),
		(drawing, 2861, 0, 4095, 0, 0),
		(drawing, 2862, 0, 4095, 0, 0),
		(drawing, 2863, 0, 4095, 0, 0),
		(drawing, 2864, 0, 4095, 0, 0),
		(drawing, 2865, 0, 4095, 0, 0),
		(drawing, 2866, 0, 4095, 0, 0),
		(drawing, 2867, 0, 4095, 0, 0),
		(drawing, 2868, 0, 4095, 0, 0),
		(drawing, 2869, 0, 4095, 0, 0),
		(drawing, 2870, 0, 4095, 0, 0),
		(drawing, 2871, 0, 4095, 0, 0),
		(drawing, 2872, 0, 4095, 0, 0),
		(drawing, 2873, 0, 4095, 0, 0),
		(drawing, 2874, 0, 4095, 0, 0),
		(drawing, 2875, 0, 4095, 0, 0),
		(drawing, 2876, 0, 4095, 0, 0),
		(drawing, 2877, 0, 4095, 0, 0),
		(drawing, 2878, 0, 4095, 0, 0),
		(drawing, 2879, 0, 4095, 0, 0),
		(drawing, 2880, 0, 4095, 0, 0),
		(drawing, 2881, 0, 4095, 0, 0),
		(drawing, 2882, 0, 4095, 0, 0),
		(drawing, 2883, 0, 4095, 0, 0),
		(drawing, 2884, 0, 4095, 0, 0),
		(drawing, 2885, 0, 4095, 0, 0),
		(drawing, 2886, 0, 4095, 0, 0),
		(drawing, 2887, 0, 4095, 0, 0),
		(drawing, 2888, 0, 4095, 0, 0),
		(drawing, 2889, 0, 4095, 0, 0),
		(drawing, 2890, 0, 4095, 0, 0),
		(drawing, 2891, 0, 4095, 0, 0),
		(drawing, 2892, 0, 4095, 0, 0),
		(drawing, 2893, 0, 4095, 0, 0),
		(drawing, 2894, 0, 4095, 0, 0),
		(drawing, 2895, 0, 4095, 0, 0),
		(drawing, 2896, 0, 4095, 0, 0),
		(drawing, 2897, 0, 4095, 0, 0),
		(drawing, 2898, 0, 4095, 0, 0),
		(drawing, 2899, 0, 4095, 0, 0),
		(drawing, 2900, 0, 4095, 0, 0),
		(drawing, 2901, 0, 4095, 0, 0),
		(drawing, 2902, 0, 4095, 0, 0),
		(drawing, 2903, 0, 4095, 0, 0),
		(drawing, 2904, 0, 4095, 0, 0),
		(drawing, 2905, 0, 4095, 0, 0),
		(drawing, 2906, 0, 4095, 0, 0),
		(drawing, 2907, 0, 4095, 0, 0),
		(drawing, 2908, 0, 4095, 0, 0),
		(drawing, 2909, 0, 4095, 0, 0),
		(drawing, 2910, 0, 4095, 0, 0),
		(drawing, 2911, 0, 4095, 0, 0),
		(drawing, 2912, 0, 4095, 0, 0),
		(drawing, 2913, 0, 4095, 0, 0),
		(drawing, 2914, 0, 4095, 0, 0),
		(drawing, 2915, 0, 4095, 0, 0),
		(drawing, 2916, 0, 4095, 0, 0),
		(drawing, 2917, 0, 4095, 0, 0),
		(drawing, 2918, 0, 4095, 0, 0),
		(drawing, 2919, 0, 4095, 0, 0),
		(drawing, 2920, 0, 4095, 0, 0),
		(drawing, 2921, 0, 4095, 0, 0),
		(drawing, 2922, 0, 4095, 0, 0),
		(drawing, 2923, 0, 4095, 0, 0),
		(drawing, 2924, 0, 4095, 0, 0),
		(drawing, 2925, 0, 4095, 0, 0),
		(drawing, 2926, 0, 4095, 0, 0),
		(drawing, 2927, 0, 4095, 0, 0),
		(drawing, 2928, 0, 4095, 0, 0),
		(drawing, 2929, 0, 4095, 0, 0),
		(drawing, 2930, 0, 4095, 0, 0),
		(drawing, 2931, 0, 4095, 0, 0),
		(drawing, 2932, 0, 4095, 0, 0),
		(drawing, 2933, 0, 4095, 0, 0),
		(drawing, 2934, 0, 4095, 0, 0),
		(drawing, 2935, 0, 4095, 0, 0),
		(drawing, 2936, 0, 4095, 0, 0),
		(drawing, 2937, 0, 4095, 0, 0),
		(drawing, 2938, 0, 4095, 0, 0),
		(drawing, 2939, 0, 4095, 0, 0),
		(drawing, 2940, 0, 4095, 0, 0),
		(drawing, 2941, 0, 4095, 0, 0),
		(drawing, 2942, 0, 4095, 0, 0),
		(drawing, 2943, 0, 4095, 0, 0),
		(drawing, 2944, 0, 4095, 0, 0),
		(drawing, 2945, 0, 4095, 0, 0),
		(drawing, 2946, 0, 4095, 0, 0),
		(drawing, 2947, 0, 4095, 0, 0),
		(drawing, 2948, 0, 4095, 0, 0),
		(drawing, 2949, 0, 4095, 0, 0),
		(drawing, 2950, 0, 4095, 0, 0),
		(drawing, 2951, 0, 4095, 0, 0),
		(drawing, 2952, 0, 4095, 0, 0),
		(drawing, 2953, 0, 4095, 0, 0),
		(drawing, 2954, 0, 4095, 0, 0),
		(drawing, 2955, 0, 4095, 0, 0),
		(drawing, 2956, 0, 4095, 0, 0),
		(drawing, 2957, 0, 4095, 0, 0),
		(drawing, 2958, 0, 4095, 0, 0),
		(drawing, 2959, 0, 4095, 0, 0),
		(drawing, 2960, 0, 4095, 0, 0),
		(drawing, 2961, 0, 4095, 0, 0),
		(drawing, 2962, 0, 4095, 0, 0),
		(drawing, 2963, 0, 4095, 0, 0),
		(drawing, 2964, 0, 4095, 0, 0),
		(drawing, 2965, 0, 4095, 0, 0),
		(drawing, 2966, 0, 4095, 0, 0),
		(drawing, 2967, 0, 4095, 0, 0),
		(drawing, 2968, 0, 4095, 0, 0),
		(drawing, 2969, 0, 4095, 0, 0),
		(drawing, 2970, 0, 4095, 0, 0),
		(drawing, 2971, 0, 4095, 0, 0),
		(drawing, 2972, 0, 4095, 0, 0),
		(drawing, 2973, 0, 4095, 0, 0),
		(drawing, 2974, 0, 4095, 0, 0),
		(drawing, 2975, 0, 4095, 0, 0),
		(drawing, 2976, 0, 4095, 0, 0),
		(drawing, 2977, 0, 4095, 0, 0),
		(drawing, 2978, 0, 4095, 0, 0),
		(drawing, 2979, 0, 4095, 0, 0),
		(drawing, 2980, 0, 4095, 0, 0),
		(drawing, 2981, 0, 4095, 0, 0),
		(drawing, 2982, 0, 4095, 0, 0),
		(drawing, 2983, 0, 4095, 0, 0),
		(drawing, 2984, 0, 4095, 0, 0),
		(drawing, 2985, 0, 4095, 0, 0),
		(drawing, 2986, 0, 4095, 0, 0),
		(drawing, 2987, 0, 4095, 0, 0),
		(drawing, 2988, 0, 4095, 0, 0),
		(drawing, 2989, 0, 4095, 0, 0),
		(drawing, 2990, 0, 4095, 0, 0),
		(drawing, 2991, 0, 4095, 0, 0),
		(drawing, 2992, 0, 4095, 0, 0),
		(drawing, 2993, 0, 4095, 0, 0),
		(drawing, 2994, 0, 4095, 0, 0),
		(drawing, 2995, 0, 4095, 0, 0),
		(drawing, 2996, 0, 4095, 0, 0),
		(drawing, 2997, 0, 4095, 0, 0),
		(drawing, 2998, 0, 4095, 0, 0),
		(drawing, 2999, 0, 4095, 0, 0),
		(drawing, 3000, 0, 4095, 0, 0),
		(drawing, 3001, 0, 4095, 0, 0),
		(drawing, 3002, 0, 4095, 0, 0),
		(drawing, 3003, 0, 4095, 0, 0),
		(drawing, 3004, 0, 4095, 0, 0),
		(drawing, 3005, 0, 4095, 0, 0),
		(drawing, 3006, 0, 4095, 0, 0),
		(drawing, 3007, 0, 4095, 0, 0),
		(drawing, 3008, 0, 4095, 0, 0),
		(drawing, 3009, 0, 4095, 0, 0),
		(drawing, 3010, 0, 4095, 0, 0),
		(drawing, 3011, 0, 4095, 0, 0),
		(drawing, 3012, 0, 4095, 0, 0),
		(drawing, 3013, 0, 4095, 0, 0),
		(drawing, 3014, 0, 4095, 0, 0),
		(drawing, 3015, 0, 4095, 0, 0),
		(drawing, 3016, 0, 4095, 0, 0),
		(drawing, 3017, 0, 4095, 0, 0),
		(drawing, 3018, 0, 4095, 0, 0),
		(drawing, 3019, 0, 4095, 0, 0),
		(drawing, 3020, 0, 4095, 0, 0),
		(drawing, 3021, 0, 4095, 0, 0),
		(drawing, 3022, 0, 4095, 0, 0),
		(drawing, 3023, 0, 4095, 0, 0),
		(drawing, 3024, 0, 4095, 0, 0),
		(drawing, 3025, 0, 4095, 0, 0),
		(drawing, 3026, 0, 4095, 0, 0),
		(drawing, 3027, 0, 4095, 0, 0),
		(drawing, 3028, 0, 4095, 0, 0),
		(drawing, 3029, 0, 4095, 0, 0),
		(drawing, 3030, 0, 4095, 0, 0),
		(drawing, 3031, 0, 4095, 0, 0),
		(drawing, 3032, 0, 4095, 0, 0),
		(drawing, 3033, 0, 4095, 0, 0),
		(drawing, 3034, 0, 4095, 0, 0),
		(drawing, 3035, 0, 4095, 0, 0),
		(drawing, 3036, 0, 4095, 0, 0),
		(drawing, 3037, 0, 4095, 0, 0),
		(drawing, 3038, 0, 4095, 0, 0),
		(drawing, 3039, 0, 4095, 0, 0),
		(drawing, 3040, 0, 4095, 0, 0),
		(drawing, 3041, 0, 4095, 0, 0),
		(drawing, 3042, 0, 4095, 0, 0),
		(drawing, 3043, 0, 4095, 0, 0),
		(drawing, 3044, 0, 4095, 0, 0),
		(drawing, 3045, 0, 4095, 0, 0),
		(drawing, 3046, 0, 4095, 0, 0),
		(drawing, 3047, 0, 4095, 0, 0),
		(drawing, 3048, 0, 4095, 0, 0),
		(drawing, 3049, 0, 4095, 0, 0),
		(drawing, 3050, 0, 4095, 0, 0),
		(drawing, 3051, 0, 4095, 0, 0),
		(drawing, 3052, 0, 4095, 0, 0),
		(drawing, 3053, 0, 4095, 0, 0),
		(drawing, 3054, 0, 4095, 0, 0),
		(drawing, 3055, 0, 4095, 0, 0),
		(drawing, 3056, 0, 4095, 0, 0),
		(drawing, 3057, 0, 4095, 0, 0),
		(drawing, 3058, 0, 4095, 0, 0),
		(drawing, 3059, 0, 4095, 0, 0),
		(drawing, 3060, 0, 4095, 0, 0),
		(drawing, 3061, 0, 4095, 0, 0),
		(drawing, 3062, 0, 4095, 0, 0),
		(drawing, 3063, 0, 4095, 0, 0),
		(drawing, 3064, 0, 4095, 0, 0),
		(drawing, 3065, 0, 4095, 0, 0),
		(drawing, 3066, 0, 4095, 0, 0),
		(drawing, 3067, 0, 4095, 0, 0),
		(drawing, 3068, 0, 4095, 0, 0),
		(drawing, 3069, 0, 4095, 0, 0),
		(drawing, 3070, 0, 4095, 0, 0),
		(drawing, 3071, 0, 4095, 0, 0),
		(drawing, 3072, 0, 4095, 0, 0),
		(drawing, 3073, 0, 4095, 0, 0),
		(drawing, 3074, 0, 4095, 0, 0),
		(drawing, 3075, 0, 4095, 0, 0),
		(drawing, 3076, 0, 4095, 0, 0),
		(drawing, 3077, 0, 4095, 0, 0),
		(drawing, 3078, 0, 4095, 0, 0),
		(drawing, 3079, 0, 4095, 0, 0),
		(drawing, 3080, 0, 4095, 0, 0),
		(drawing, 3081, 0, 4095, 0, 0),
		(drawing, 3082, 0, 4095, 0, 0),
		(drawing, 3083, 0, 4095, 0, 0),
		(drawing, 3084, 0, 4095, 0, 0),
		(drawing, 3085, 0, 4095, 0, 0),
		(drawing, 3086, 0, 4095, 0, 0),
		(drawing, 3087, 0, 4095, 0, 0),
		(drawing, 3088, 0, 4095, 0, 0),
		(drawing, 3089, 0, 4095, 0, 0),
		(drawing, 3090, 0, 4095, 0, 0),
		(drawing, 3091, 0, 4095, 0, 0),
		(drawing, 3092, 0, 4095, 0, 0),
		(drawing, 3093, 0, 4095, 0, 0),
		(drawing, 3094, 0, 4095, 0, 0),
		(drawing, 3095, 0, 4095, 0, 0),
		(drawing, 3096, 0, 4095, 0, 0),
		(drawing, 3097, 0, 4095, 0, 0),
		(drawing, 3098, 0, 4095, 0, 0),
		(drawing, 3099, 0, 4095, 0, 0),
		(drawing, 3100, 0, 4095, 0, 0),
		(drawing, 3101, 0, 4095, 0, 0),
		(drawing, 3102, 0, 4095, 0, 0),
		(drawing, 3103, 0, 4095, 0, 0),
		(drawing, 3104, 0, 4095, 0, 0),
		(drawing, 3105, 0, 4095, 0, 0),
		(drawing, 3106, 0, 4095, 0, 0),
		(drawing, 3107, 0, 4095, 0, 0),
		(drawing, 3108, 0, 4095, 0, 0),
		(drawing, 3109, 0, 4095, 0, 0),
		(drawing, 3110, 0, 4095, 0, 0),
		(drawing, 3111, 0, 4095, 0, 0),
		(drawing, 3112, 0, 4095, 0, 0),
		(drawing, 3113, 0, 4095, 0, 0),
		(drawing, 3114, 0, 4095, 0, 0),
		(drawing, 3115, 0, 4095, 0, 0),
		(drawing, 3116, 0, 4095, 0, 0),
		(drawing, 3117, 0, 4095, 0, 0),
		(drawing, 3118, 0, 4095, 0, 0),
		(drawing, 3119, 0, 4095, 0, 0),
		(drawing, 3120, 0, 4095, 0, 0),
		(drawing, 3121, 0, 4095, 0, 0),
		(drawing, 3122, 0, 4095, 0, 0),
		(drawing, 3123, 0, 4095, 0, 0),
		(drawing, 3124, 0, 4095, 0, 0),
		(drawing, 3125, 0, 4095, 0, 0),
		(drawing, 3126, 0, 4095, 0, 0),
		(drawing, 3127, 0, 4095, 0, 0),
		(drawing, 3128, 0, 4095, 0, 0),
		(drawing, 3129, 0, 4095, 0, 0),
		(drawing, 3130, 0, 4095, 0, 0),
		(drawing, 3131, 0, 4095, 0, 0),
		(drawing, 3132, 0, 4095, 0, 0),
		(drawing, 3133, 0, 4095, 0, 0),
		(drawing, 3134, 0, 4095, 0, 0),
		(drawing, 3135, 0, 4095, 0, 0),
		(drawing, 3136, 0, 4095, 0, 0),
		(drawing, 3137, 0, 4095, 0, 0),
		(drawing, 3138, 0, 4095, 0, 0),
		(drawing, 3139, 0, 4095, 0, 0),
		(drawing, 3140, 0, 4095, 0, 0),
		(drawing, 3141, 0, 4095, 0, 0),
		(drawing, 3142, 0, 4095, 0, 0),
		(drawing, 3143, 0, 4095, 0, 0),
		(drawing, 3144, 0, 4095, 0, 0),
		(drawing, 3145, 0, 4095, 0, 0),
		(drawing, 3146, 0, 4095, 0, 0),
		(drawing, 3147, 0, 4095, 0, 0),
		(drawing, 3148, 0, 4095, 0, 0),
		(drawing, 3149, 0, 4095, 0, 0),
		(drawing, 3150, 0, 4095, 0, 0),
		(drawing, 3151, 0, 4095, 0, 0),
		(drawing, 3152, 0, 4095, 0, 0),
		(drawing, 3153, 0, 4095, 0, 0),
		(drawing, 3154, 0, 4095, 0, 0),
		(drawing, 3155, 0, 4095, 0, 0),
		(drawing, 3156, 0, 4095, 0, 0),
		(drawing, 3157, 0, 4095, 0, 0),
		(drawing, 3158, 0, 4095, 0, 0),
		(drawing, 3159, 0, 4095, 0, 0),
		(drawing, 3160, 0, 4095, 0, 0),
		(drawing, 3161, 0, 4095, 0, 0),
		(drawing, 3162, 0, 4095, 0, 0),
		(drawing, 3163, 0, 4095, 0, 0),
		(drawing, 3164, 0, 4095, 0, 0),
		(drawing, 3165, 0, 4095, 0, 0),
		(drawing, 3166, 0, 4095, 0, 0),
		(drawing, 3167, 0, 4095, 0, 0),
		(drawing, 3168, 0, 4095, 0, 0),
		(drawing, 3169, 0, 4095, 0, 0),
		(drawing, 3170, 0, 4095, 0, 0),
		(drawing, 3171, 0, 4095, 0, 0),
		(drawing, 3172, 0, 4095, 0, 0),
		(drawing, 3173, 0, 4095, 0, 0),
		(drawing, 3174, 0, 4095, 0, 0),
		(drawing, 3175, 0, 4095, 0, 0),
		(drawing, 3176, 0, 4095, 0, 0),
		(drawing, 3177, 0, 4095, 0, 0),
		(drawing, 3178, 0, 4095, 0, 0),
		(drawing, 3179, 0, 4095, 0, 0),
		(drawing, 3180, 0, 4095, 0, 0),
		(drawing, 3181, 0, 4095, 0, 0),
		(drawing, 3182, 0, 4095, 0, 0),
		(drawing, 3183, 0, 4095, 0, 0),
		(drawing, 3184, 0, 4095, 0, 0),
		(drawing, 3185, 0, 4095, 0, 0),
		(drawing, 3186, 0, 4095, 0, 0),
		(drawing, 3187, 0, 4095, 0, 0),
		(drawing, 3188, 0, 4095, 0, 0),
		(drawing, 3189, 0, 4095, 0, 0),
		(drawing, 3190, 0, 4095, 0, 0),
		(drawing, 3191, 0, 4095, 0, 0),
		(drawing, 3192, 0, 4095, 0, 0),
		(drawing, 3193, 0, 4095, 0, 0),
		(drawing, 3194, 0, 4095, 0, 0),
		(drawing, 3195, 0, 4095, 0, 0),
		(drawing, 3196, 0, 4095, 0, 0),
		(drawing, 3197, 0, 4095, 0, 0),
		(drawing, 3198, 0, 4095, 0, 0),
		(drawing, 3199, 0, 4095, 0, 0),
		(drawing, 3200, 0, 4095, 0, 0),
		(drawing, 3201, 0, 4095, 0, 0),
		(drawing, 3202, 0, 4095, 0, 0),
		(drawing, 3203, 0, 4095, 0, 0),
		(drawing, 3204, 0, 4095, 0, 0),
		(drawing, 3205, 0, 4095, 0, 0),
		(drawing, 3206, 0, 4095, 0, 0),
		(drawing, 3207, 0, 4095, 0, 0),
		(drawing, 3208, 0, 4095, 0, 0),
		(drawing, 3209, 0, 4095, 0, 0),
		(drawing, 3210, 0, 4095, 0, 0),
		(drawing, 3211, 0, 4095, 0, 0),
		(drawing, 3212, 0, 4095, 0, 0),
		(drawing, 3213, 0, 4095, 0, 0),
		(drawing, 3214, 0, 4095, 0, 0),
		(drawing, 3215, 0, 4095, 0, 0),
		(drawing, 3216, 0, 4095, 0, 0),
		(drawing, 3217, 0, 4095, 0, 0),
		(drawing, 3218, 0, 4095, 0, 0),
		(drawing, 3219, 0, 4095, 0, 0),
		(drawing, 3220, 0, 4095, 0, 0),
		(drawing, 3221, 0, 4095, 0, 0),
		(drawing, 3222, 0, 4095, 0, 0),
		(drawing, 3223, 0, 4095, 0, 0),
		(drawing, 3224, 0, 4095, 0, 0),
		(drawing, 3225, 0, 4095, 0, 0),
		(drawing, 3226, 0, 4095, 0, 0),
		(drawing, 3227, 0, 4095, 0, 0),
		(drawing, 3228, 0, 4095, 0, 0),
		(drawing, 3229, 0, 4095, 0, 0),
		(drawing, 3230, 0, 4095, 0, 0),
		(drawing, 3231, 0, 4095, 0, 0),
		(drawing, 3232, 0, 4095, 0, 0),
		(drawing, 3233, 0, 4095, 0, 0),
		(drawing, 3234, 0, 4095, 0, 0),
		(drawing, 3235, 0, 4095, 0, 0),
		(drawing, 3236, 0, 4095, 0, 0),
		(drawing, 3237, 0, 4095, 0, 0),
		(drawing, 3238, 0, 4095, 0, 0),
		(drawing, 3239, 0, 4095, 0, 0),
		(drawing, 3240, 0, 4095, 0, 0),
		(drawing, 3241, 0, 4095, 0, 0),
		(drawing, 3242, 0, 4095, 0, 0),
		(drawing, 3243, 0, 4095, 0, 0),
		(drawing, 3244, 0, 4095, 0, 0),
		(drawing, 3245, 0, 4095, 0, 0),
		(drawing, 3246, 0, 4095, 0, 0),
		(drawing, 3247, 0, 4095, 0, 0),
		(drawing, 3248, 0, 4095, 0, 0),
		(drawing, 3249, 0, 4095, 0, 0),
		(drawing, 3250, 0, 4095, 0, 0),
		(drawing, 3251, 0, 4095, 0, 0),
		(drawing, 3252, 0, 4095, 0, 0),
		(drawing, 3253, 0, 4095, 0, 0),
		(drawing, 3254, 0, 4095, 0, 0),
		(drawing, 3255, 0, 4095, 0, 0),
		(drawing, 3256, 0, 4095, 0, 0),
		(drawing, 3257, 0, 4095, 0, 0),
		(drawing, 3258, 0, 4095, 0, 0),
		(drawing, 3259, 0, 4095, 0, 0),
		(drawing, 3260, 0, 4095, 0, 0),
		(drawing, 3261, 0, 4095, 0, 0),
		(drawing, 3262, 0, 4095, 0, 0),
		(drawing, 3263, 0, 4095, 0, 0),
		(drawing, 3264, 0, 4095, 0, 0),
		(drawing, 3265, 0, 4095, 0, 0),
		(drawing, 3266, 0, 4095, 0, 0),
		(drawing, 3267, 0, 4095, 0, 0),
		(drawing, 3268, 0, 4095, 0, 0),
		(drawing, 3269, 0, 4095, 0, 0),
		(drawing, 3270, 0, 4095, 0, 0),
		(drawing, 3271, 0, 4095, 0, 0),
		(drawing, 3272, 0, 4095, 0, 0),
		(drawing, 3273, 0, 4095, 0, 0),
		(drawing, 3274, 0, 4095, 0, 0),
		(drawing, 3275, 0, 4095, 0, 0),
		(drawing, 3276, 0, 4095, 0, 0),
		(drawing, 3277, 0, 4095, 0, 0),
		(drawing, 3278, 0, 4095, 0, 0),
		(drawing, 3279, 0, 4095, 0, 0),
		(drawing, 3280, 0, 4095, 0, 0),
		(drawing, 3281, 0, 4095, 0, 0),
		(drawing, 3282, 0, 4095, 0, 0),
		(drawing, 3283, 0, 4095, 0, 0),
		(drawing, 3284, 0, 4095, 0, 0),
		(drawing, 3285, 0, 4095, 0, 0),
		(drawing, 3286, 0, 4095, 0, 0),
		(drawing, 3287, 0, 4095, 0, 0),
		(drawing, 3288, 0, 4095, 0, 0),
		(drawing, 3289, 0, 4095, 0, 0),
		(drawing, 3290, 0, 4095, 0, 0),
		(drawing, 3291, 0, 4095, 0, 0),
		(drawing, 3292, 0, 4095, 0, 0),
		(drawing, 3293, 0, 4095, 0, 0),
		(drawing, 3294, 0, 4095, 0, 0),
		(drawing, 3295, 0, 4095, 0, 0),
		(drawing, 3296, 0, 4095, 0, 0),
		(drawing, 3297, 0, 4095, 0, 0),
		(drawing, 3298, 0, 4095, 0, 0),
		(drawing, 3299, 0, 4095, 0, 0),
		(drawing, 3300, 0, 4095, 0, 0),
		(drawing, 3301, 0, 4095, 0, 0),
		(drawing, 3302, 0, 4095, 0, 0),
		(drawing, 3303, 0, 4095, 0, 0),
		(drawing, 3304, 0, 4095, 0, 0),
		(drawing, 3305, 0, 4095, 0, 0),
		(drawing, 3306, 0, 4095, 0, 0),
		(drawing, 3307, 0, 4095, 0, 0),
		(drawing, 3308, 0, 4095, 0, 0),
		(drawing, 3309, 0, 4095, 0, 0),
		(drawing, 3310, 0, 4095, 0, 0),
		(drawing, 3311, 0, 4095, 0, 0),
		(drawing, 3312, 0, 4095, 0, 0),
		(drawing, 3313, 0, 4095, 0, 0),
		(drawing, 3314, 0, 4095, 0, 0),
		(drawing, 3315, 0, 4095, 0, 0),
		(drawing, 3316, 0, 4095, 0, 0),
		(drawing, 3317, 0, 4095, 0, 0),
		(drawing, 3318, 0, 4095, 0, 0),
		(drawing, 3319, 0, 4095, 0, 0),
		(drawing, 3320, 0, 4095, 0, 0),
		(drawing, 3321, 0, 4095, 0, 0),
		(drawing, 3322, 0, 4095, 0, 0),
		(drawing, 3323, 0, 4095, 0, 0),
		(drawing, 3324, 0, 4095, 0, 0),
		(drawing, 3325, 0, 4095, 0, 0),
		(drawing, 3326, 0, 4095, 0, 0),
		(drawing, 3327, 0, 4095, 0, 0),
		(drawing, 3328, 0, 4095, 0, 0),
		(drawing, 3329, 0, 4095, 0, 0),
		(drawing, 3330, 0, 4095, 0, 0),
		(drawing, 3331, 0, 4095, 0, 0),
		(drawing, 3332, 0, 4095, 0, 0),
		(drawing, 3333, 0, 4095, 0, 0),
		(drawing, 3334, 0, 4095, 0, 0),
		(drawing, 3335, 0, 4095, 0, 0),
		(drawing, 3336, 0, 4095, 0, 0),
		(drawing, 3337, 0, 4095, 0, 0),
		(drawing, 3338, 0, 4095, 0, 0),
		(drawing, 3339, 0, 4095, 0, 0),
		(drawing, 3340, 0, 4095, 0, 0),
		(drawing, 3341, 0, 4095, 0, 0),
		(drawing, 3342, 0, 4095, 0, 0),
		(drawing, 3343, 0, 4095, 0, 0),
		(drawing, 3344, 0, 4095, 0, 0),
		(drawing, 3345, 0, 4095, 0, 0),
		(drawing, 3346, 0, 4095, 0, 0),
		(drawing, 3347, 0, 4095, 0, 0),
		(drawing, 3348, 0, 4095, 0, 0),
		(drawing, 3349, 0, 4095, 0, 0),
		(drawing, 3350, 0, 4095, 0, 0),
		(drawing, 3351, 0, 4095, 0, 0),
		(drawing, 3352, 0, 4095, 0, 0),
		(drawing, 3353, 0, 4095, 0, 0),
		(drawing, 3354, 0, 4095, 0, 0),
		(drawing, 3355, 0, 4095, 0, 0),
		(drawing, 3356, 0, 4095, 0, 0),
		(drawing, 3357, 0, 4095, 0, 0),
		(drawing, 3358, 0, 4095, 0, 0),
		(drawing, 3359, 0, 4095, 0, 0),
		(drawing, 3360, 0, 4095, 0, 0),
		(drawing, 3361, 0, 4095, 0, 0),
		(drawing, 3362, 0, 4095, 0, 0),
		(drawing, 3363, 0, 4095, 0, 0),
		(drawing, 3364, 0, 4095, 0, 0),
		(drawing, 3365, 0, 4095, 0, 0),
		(drawing, 3366, 0, 4095, 0, 0),
		(drawing, 3367, 0, 4095, 0, 0),
		(drawing, 3368, 0, 4095, 0, 0),
		(drawing, 3369, 0, 4095, 0, 0),
		(drawing, 3370, 0, 4095, 0, 0),
		(drawing, 3371, 0, 4095, 0, 0),
		(drawing, 3372, 0, 4095, 0, 0),
		(drawing, 3373, 0, 4095, 0, 0),
		(drawing, 3374, 0, 4095, 0, 0),
		(drawing, 3375, 0, 4095, 0, 0),
		(drawing, 3376, 0, 4095, 0, 0),
		(drawing, 3377, 0, 4095, 0, 0),
		(drawing, 3378, 0, 4095, 0, 0),
		(drawing, 3379, 0, 4095, 0, 0),
		(drawing, 3380, 0, 4095, 0, 0),
		(drawing, 3381, 0, 4095, 0, 0),
		(drawing, 3382, 0, 4095, 0, 0),
		(drawing, 3383, 0, 4095, 0, 0),
		(drawing, 3384, 0, 4095, 0, 0),
		(drawing, 3385, 0, 4095, 0, 0),
		(drawing, 3386, 0, 4095, 0, 0),
		(drawing, 3387, 0, 4095, 0, 0),
		(drawing, 3388, 0, 4095, 0, 0),
		(drawing, 3389, 0, 4095, 0, 0),
		(drawing, 3390, 0, 4095, 0, 0),
		(drawing, 3391, 0, 4095, 0, 0),
		(drawing, 3392, 0, 4095, 0, 0),
		(drawing, 3393, 0, 4095, 0, 0),
		(drawing, 3394, 0, 4095, 0, 0),
		(drawing, 3395, 0, 4095, 0, 0),
		(drawing, 3396, 0, 4095, 0, 0),
		(drawing, 3397, 0, 4095, 0, 0),
		(drawing, 3398, 0, 4095, 0, 0),
		(drawing, 3399, 0, 4095, 0, 0),
		(drawing, 3400, 0, 4095, 0, 0),
		(drawing, 3401, 0, 4095, 0, 0),
		(drawing, 3402, 0, 4095, 0, 0),
		(drawing, 3403, 0, 4095, 0, 0),
		(drawing, 3404, 0, 4095, 0, 0),
		(drawing, 3405, 0, 4095, 0, 0),
		(drawing, 3406, 0, 4095, 0, 0),
		(drawing, 3407, 0, 4095, 0, 0),
		(drawing, 3408, 0, 4095, 0, 0),
		(drawing, 3409, 0, 4095, 0, 0),
		(drawing, 3410, 0, 4095, 0, 0),
		(drawing, 3411, 0, 4095, 0, 0),
		(drawing, 3412, 0, 4095, 0, 0),
		(drawing, 3413, 0, 4095, 0, 0),
		(drawing, 3414, 0, 4095, 0, 0),
		(drawing, 3415, 0, 4095, 0, 0),
		(drawing, 3416, 0, 4095, 0, 0),
		(drawing, 3417, 0, 4095, 0, 0),
		(drawing, 3418, 0, 4095, 0, 0),
		(drawing, 3419, 0, 4095, 0, 0),
		(drawing, 3420, 0, 4095, 0, 0),
		(drawing, 3421, 0, 4095, 0, 0),
		(drawing, 3422, 0, 4095, 0, 0),
		(drawing, 3423, 0, 4095, 0, 0),
		(drawing, 3424, 0, 4095, 0, 0),
		(drawing, 3425, 0, 4095, 0, 0),
		(drawing, 3426, 0, 4095, 0, 0),
		(drawing, 3427, 0, 4095, 0, 0),
		(drawing, 3428, 0, 4095, 0, 0),
		(drawing, 3429, 0, 4095, 0, 0),
		(drawing, 3430, 0, 4095, 0, 0),
		(drawing, 3431, 0, 4095, 0, 0),
		(drawing, 3432, 0, 4095, 0, 0),
		(drawing, 3433, 0, 4095, 0, 0),
		(drawing, 3434, 0, 4095, 0, 0),
		(drawing, 3435, 0, 4095, 0, 0),
		(drawing, 3436, 0, 4095, 0, 0),
		(drawing, 3437, 0, 4095, 0, 0),
		(drawing, 3438, 0, 4095, 0, 0),
		(drawing, 3439, 0, 4095, 0, 0),
		(drawing, 3440, 0, 4095, 0, 0),
		(drawing, 3441, 0, 4095, 0, 0),
		(drawing, 3442, 0, 4095, 0, 0),
		(drawing, 3443, 0, 4095, 0, 0),
		(drawing, 3444, 0, 4095, 0, 0),
		(drawing, 3445, 0, 4095, 0, 0),
		(drawing, 3446, 0, 4095, 0, 0),
		(drawing, 3447, 0, 4095, 0, 0),
		(drawing, 3448, 0, 4095, 0, 0),
		(drawing, 3449, 0, 4095, 0, 0),
		(drawing, 3450, 0, 4095, 0, 0),
		(drawing, 3451, 0, 4095, 0, 0),
		(drawing, 3452, 0, 4095, 0, 0),
		(drawing, 3453, 0, 4095, 0, 0),
		(drawing, 3454, 0, 4095, 0, 0),
		(drawing, 3455, 0, 4095, 0, 0),
		(drawing, 3456, 0, 4095, 0, 0),
		(drawing, 3457, 0, 4095, 0, 0),
		(drawing, 3458, 0, 4095, 0, 0),
		(drawing, 3459, 0, 4095, 0, 0),
		(drawing, 3460, 0, 4095, 0, 0),
		(drawing, 3461, 0, 4095, 0, 0),
		(drawing, 3462, 0, 4095, 0, 0),
		(drawing, 3463, 0, 4095, 0, 0),
		(drawing, 3464, 0, 4095, 0, 0),
		(drawing, 3465, 0, 4095, 0, 0),
		(drawing, 3466, 0, 4095, 0, 0),
		(drawing, 3467, 0, 4095, 0, 0),
		(drawing, 3468, 0, 4095, 0, 0),
		(drawing, 3469, 0, 4095, 0, 0),
		(drawing, 3470, 0, 4095, 0, 0),
		(drawing, 3471, 0, 4095, 0, 0),
		(drawing, 3472, 0, 4095, 0, 0),
		(drawing, 3473, 0, 4095, 0, 0),
		(drawing, 3474, 0, 4095, 0, 0),
		(drawing, 3475, 0, 4095, 0, 0),
		(drawing, 3476, 0, 4095, 0, 0),
		(drawing, 3477, 0, 4095, 0, 0),
		(drawing, 3478, 0, 4095, 0, 0),
		(drawing, 3479, 0, 4095, 0, 0),
		(drawing, 3480, 0, 4095, 0, 0),
		(drawing, 3481, 0, 4095, 0, 0),
		(drawing, 3482, 0, 4095, 0, 0),
		(drawing, 3483, 0, 4095, 0, 0),
		(drawing, 3484, 0, 4095, 0, 0),
		(drawing, 3485, 0, 4095, 0, 0),
		(drawing, 3486, 0, 4095, 0, 0),
		(drawing, 3487, 0, 4095, 0, 0),
		(drawing, 3488, 0, 4095, 0, 0),
		(drawing, 3489, 0, 4095, 0, 0),
		(drawing, 3490, 0, 4095, 0, 0),
		(drawing, 3491, 0, 4095, 0, 0),
		(drawing, 3492, 0, 4095, 0, 0),
		(drawing, 3493, 0, 4095, 0, 0),
		(drawing, 3494, 0, 4095, 0, 0),
		(drawing, 3495, 0, 4095, 0, 0),
		(drawing, 3496, 0, 4095, 0, 0),
		(drawing, 3497, 0, 4095, 0, 0),
		(drawing, 3498, 0, 4095, 0, 0),
		(drawing, 3499, 0, 4095, 0, 0),
		(drawing, 3500, 0, 4095, 0, 0),
		(drawing, 3501, 0, 4095, 0, 0),
		(drawing, 3502, 0, 4095, 0, 0),
		(drawing, 3503, 0, 4095, 0, 0),
		(drawing, 3504, 0, 4095, 0, 0),
		(drawing, 3505, 0, 4095, 0, 0),
		(drawing, 3506, 0, 4095, 0, 0),
		(drawing, 3507, 0, 4095, 0, 0),
		(drawing, 3508, 0, 4095, 0, 0),
		(drawing, 3509, 0, 4095, 0, 0),
		(drawing, 3510, 0, 4095, 0, 0),
		(drawing, 3511, 0, 4095, 0, 0),
		(drawing, 3512, 0, 4095, 0, 0),
		(drawing, 3513, 0, 4095, 0, 0),
		(drawing, 3514, 0, 4095, 0, 0),
		(drawing, 3515, 0, 4095, 0, 0),
		(drawing, 3516, 0, 4095, 0, 0),
		(drawing, 3517, 0, 4095, 0, 0),
		(drawing, 3518, 0, 4095, 0, 0),
		(drawing, 3519, 0, 4095, 0, 0),
		(drawing, 3520, 0, 4095, 0, 0),
		(drawing, 3521, 0, 4095, 0, 0),
		(drawing, 3522, 0, 4095, 0, 0),
		(drawing, 3523, 0, 4095, 0, 0),
		(drawing, 3524, 0, 4095, 0, 0),
		(drawing, 3525, 0, 4095, 0, 0),
		(drawing, 3526, 0, 4095, 0, 0),
		(drawing, 3527, 0, 4095, 0, 0),
		(drawing, 3528, 0, 4095, 0, 0),
		(drawing, 3529, 0, 4095, 0, 0),
		(drawing, 3530, 0, 4095, 0, 0),
		(drawing, 3531, 0, 4095, 0, 0),
		(drawing, 3532, 0, 4095, 0, 0),
		(drawing, 3533, 0, 4095, 0, 0),
		(drawing, 3534, 0, 4095, 0, 0),
		(drawing, 3535, 0, 4095, 0, 0),
		(drawing, 3536, 0, 4095, 0, 0),
		(drawing, 3537, 0, 4095, 0, 0),
		(drawing, 3538, 0, 4095, 0, 0),
		(drawing, 3539, 0, 4095, 0, 0),
		(drawing, 3540, 0, 4095, 0, 0),
		(drawing, 3541, 0, 4095, 0, 0),
		(drawing, 3542, 0, 4095, 0, 0),
		(drawing, 3543, 0, 4095, 0, 0),
		(drawing, 3544, 0, 4095, 0, 0),
		(drawing, 3545, 0, 4095, 0, 0),
		(drawing, 3546, 0, 4095, 0, 0),
		(drawing, 3547, 0, 4095, 0, 0),
		(drawing, 3548, 0, 4095, 0, 0),
		(drawing, 3549, 0, 4095, 0, 0),
		(drawing, 3550, 0, 4095, 0, 0),
		(drawing, 3551, 0, 4095, 0, 0),
		(drawing, 3552, 0, 4095, 0, 0),
		(drawing, 3553, 0, 4095, 0, 0),
		(drawing, 3554, 0, 4095, 0, 0),
		(drawing, 3555, 0, 4095, 0, 0),
		(drawing, 3556, 0, 4095, 0, 0),
		(drawing, 3557, 0, 4095, 0, 0),
		(drawing, 3558, 0, 4095, 0, 0),
		(drawing, 3559, 0, 4095, 0, 0),
		(drawing, 3560, 0, 4095, 0, 0),
		(drawing, 3561, 0, 4095, 0, 0),
		(drawing, 3562, 0, 4095, 0, 0),
		(drawing, 3563, 0, 4095, 0, 0),
		(drawing, 3564, 0, 4095, 0, 0),
		(drawing, 3565, 0, 4095, 0, 0),
		(drawing, 3566, 0, 4095, 0, 0),
		(drawing, 3567, 0, 4095, 0, 0),
		(drawing, 3568, 0, 4095, 0, 0),
		(drawing, 3569, 0, 4095, 0, 0),
		(drawing, 3570, 0, 4095, 0, 0),
		(drawing, 3571, 0, 4095, 0, 0),
		(drawing, 3572, 0, 4095, 0, 0),
		(drawing, 3573, 0, 4095, 0, 0),
		(drawing, 3574, 0, 4095, 0, 0),
		(drawing, 3575, 0, 4095, 0, 0),
		(drawing, 3576, 0, 4095, 0, 0),
		(drawing, 3577, 0, 4095, 0, 0),
		(drawing, 3578, 0, 4095, 0, 0),
		(drawing, 3579, 0, 4095, 0, 0),
		(drawing, 3580, 0, 4095, 0, 0),
		(drawing, 3581, 0, 4095, 0, 0),
		(drawing, 3582, 0, 4095, 0, 0),
		(drawing, 3583, 0, 4095, 0, 0),
		(drawing, 3584, 0, 4095, 0, 0),
		(drawing, 3585, 0, 4095, 0, 0),
		(drawing, 3586, 0, 4095, 0, 0),
		(drawing, 3587, 0, 4095, 0, 0),
		(drawing, 3588, 0, 4095, 0, 0),
		(drawing, 3589, 0, 4095, 0, 0),
		(drawing, 3590, 0, 4095, 0, 0),
		(drawing, 3591, 0, 4095, 0, 0),
		(drawing, 3592, 0, 4095, 0, 0),
		(drawing, 3593, 0, 4095, 0, 0),
		(drawing, 3594, 0, 4095, 0, 0),
		(drawing, 3595, 0, 4095, 0, 0),
		(drawing, 3596, 0, 4095, 0, 0),
		(drawing, 3597, 0, 4095, 0, 0),
		(drawing, 3598, 0, 4095, 0, 0),
		(drawing, 3599, 0, 4095, 0, 0),
		(drawing, 3600, 0, 4095, 0, 0),
		(drawing, 3601, 0, 4095, 0, 0),
		(drawing, 3602, 0, 4095, 0, 0),
		(drawing, 3603, 0, 4095, 0, 0),
		(drawing, 3604, 0, 4095, 0, 0),
		(drawing, 3605, 0, 4095, 0, 0),
		(drawing, 3606, 0, 4095, 0, 0),
		(drawing, 3607, 0, 4095, 0, 0),
		(drawing, 3608, 0, 4095, 0, 0),
		(drawing, 3609, 0, 4095, 0, 0),
		(drawing, 3610, 0, 4095, 0, 0),
		(drawing, 3611, 0, 4095, 0, 0),
		(drawing, 3612, 0, 4095, 0, 0),
		(drawing, 3613, 0, 4095, 0, 0),
		(drawing, 3614, 0, 4095, 0, 0),
		(drawing, 3615, 0, 4095, 0, 0),
		(drawing, 3616, 0, 4095, 0, 0),
		(drawing, 3617, 0, 4095, 0, 0),
		(drawing, 3618, 0, 4095, 0, 0),
		(drawing, 3619, 0, 4095, 0, 0),
		(drawing, 3620, 0, 4095, 0, 0),
		(drawing, 3621, 0, 4095, 0, 0),
		(drawing, 3622, 0, 4095, 0, 0),
		(drawing, 3623, 0, 4095, 0, 0),
		(drawing, 3624, 0, 4095, 0, 0),
		(drawing, 3625, 0, 4095, 0, 0),
		(drawing, 3626, 0, 4095, 0, 0),
		(drawing, 3627, 0, 4095, 0, 0),
		(drawing, 3628, 0, 4095, 0, 0),
		(drawing, 3629, 0, 4095, 0, 0),
		(drawing, 3630, 0, 4095, 0, 0),
		(drawing, 3631, 0, 4095, 0, 0),
		(drawing, 3632, 0, 4095, 0, 0),
		(drawing, 3633, 0, 4095, 0, 0),
		(drawing, 3634, 0, 4095, 0, 0),
		(drawing, 3635, 0, 4095, 0, 0),
		(drawing, 3636, 0, 4095, 0, 0),
		(drawing, 3637, 0, 4095, 0, 0),
		(drawing, 3638, 0, 4095, 0, 0),
		(drawing, 3639, 0, 4095, 0, 0),
		(drawing, 3640, 0, 4095, 0, 0),
		(drawing, 3641, 0, 4095, 0, 0),
		(drawing, 3642, 0, 4095, 0, 0),
		(drawing, 3643, 0, 4095, 0, 0),
		(drawing, 3644, 0, 4095, 0, 0),
		(drawing, 3645, 0, 4095, 0, 0),
		(drawing, 3646, 0, 4095, 0, 0),
		(drawing, 3647, 0, 4095, 0, 0),
		(drawing, 3648, 0, 4095, 0, 0),
		(drawing, 3649, 0, 4095, 0, 0),
		(drawing, 3650, 0, 4095, 0, 0),
		(drawing, 3651, 0, 4095, 0, 0),
		(drawing, 3652, 0, 4095, 0, 0),
		(drawing, 3653, 0, 4095, 0, 0),
		(drawing, 3654, 0, 4095, 0, 0),
		(drawing, 3655, 0, 4095, 0, 0),
		(drawing, 3656, 0, 4095, 0, 0),
		(drawing, 3657, 0, 4095, 0, 0),
		(drawing, 3658, 0, 4095, 0, 0),
		(drawing, 3659, 0, 4095, 0, 0),
		(drawing, 3660, 0, 4095, 0, 0),
		(drawing, 3661, 0, 4095, 0, 0),
		(drawing, 3662, 0, 4095, 0, 0),
		(drawing, 3663, 0, 4095, 0, 0),
		(drawing, 3664, 0, 4095, 0, 0),
		(drawing, 3665, 0, 4095, 0, 0),
		(drawing, 3666, 0, 4095, 0, 0),
		(drawing, 3667, 0, 4095, 0, 0),
		(drawing, 3668, 0, 4095, 0, 0),
		(drawing, 3669, 0, 4095, 0, 0),
		(drawing, 3670, 0, 4095, 0, 0),
		(drawing, 3671, 0, 4095, 0, 0),
		(drawing, 3672, 0, 4095, 0, 0),
		(drawing, 3673, 0, 4095, 0, 0),
		(drawing, 3674, 0, 4095, 0, 0),
		(drawing, 3675, 0, 4095, 0, 0),
		(drawing, 3676, 0, 4095, 0, 0),
		(drawing, 3677, 0, 4095, 0, 0),
		(drawing, 3678, 0, 4095, 0, 0),
		(drawing, 3679, 0, 4095, 0, 0),
		(drawing, 3680, 0, 4095, 0, 0),
		(drawing, 3681, 0, 4095, 0, 0),
		(drawing, 3682, 0, 4095, 0, 0),
		(drawing, 3683, 0, 4095, 0, 0),
		(drawing, 3684, 0, 4095, 0, 0),
		(drawing, 3685, 0, 4095, 0, 0),
		(drawing, 3686, 0, 4095, 0, 0),
		(drawing, 3687, 0, 4095, 0, 0),
		(drawing, 3688, 0, 4095, 0, 0),
		(drawing, 3689, 0, 4095, 0, 0),
		(drawing, 3690, 0, 4095, 0, 0),
		(drawing, 3691, 0, 4095, 0, 0),
		(drawing, 3692, 0, 4095, 0, 0),
		(drawing, 3693, 0, 4095, 0, 0),
		(drawing, 3694, 0, 4095, 0, 0),
		(drawing, 3695, 0, 4095, 0, 0),
		(drawing, 3696, 0, 4095, 0, 0),
		(drawing, 3697, 0, 4095, 0, 0),
		(drawing, 3698, 0, 4095, 0, 0),
		(drawing, 3699, 0, 4095, 0, 0),
		(drawing, 3700, 0, 4095, 0, 0),
		(drawing, 3701, 0, 4095, 0, 0),
		(drawing, 3702, 0, 4095, 0, 0),
		(drawing, 3703, 0, 4095, 0, 0),
		(drawing, 3704, 0, 4095, 0, 0),
		(drawing, 3705, 0, 4095, 0, 0),
		(drawing, 3706, 0, 4095, 0, 0),
		(drawing, 3707, 0, 4095, 0, 0),
		(drawing, 3708, 0, 4095, 0, 0),
		(drawing, 3709, 0, 4095, 0, 0),
		(drawing, 3710, 0, 4095, 0, 0),
		(drawing, 3711, 0, 4095, 0, 0),
		(drawing, 3712, 0, 4095, 0, 0),
		(drawing, 3713, 0, 4095, 0, 0),
		(drawing, 3714, 0, 4095, 0, 0),
		(drawing, 3715, 0, 4095, 0, 0),
		(drawing, 3716, 0, 4095, 0, 0),
		(drawing, 3717, 0, 4095, 0, 0),
		(drawing, 3718, 0, 4095, 0, 0),
		(drawing, 3719, 0, 4095, 0, 0),
		(drawing, 3720, 0, 4095, 0, 0),
		(drawing, 3721, 0, 4095, 0, 0),
		(drawing, 3722, 0, 4095, 0, 0),
		(drawing, 3723, 0, 4095, 0, 0),
		(drawing, 3724, 0, 4095, 0, 0),
		(drawing, 3725, 0, 4095, 0, 0),
		(drawing, 3726, 0, 4095, 0, 0),
		(drawing, 3727, 0, 4095, 0, 0),
		(drawing, 3728, 0, 4095, 0, 0),
		(drawing, 3729, 0, 4095, 0, 0),
		(drawing, 3730, 0, 4095, 0, 0),
		(drawing, 3731, 0, 4095, 0, 0),
		(drawing, 3732, 0, 4095, 0, 0),
		(drawing, 3733, 0, 4095, 0, 0),
		(drawing, 3734, 0, 4095, 0, 0),
		(drawing, 3735, 0, 4095, 0, 0),
		(drawing, 3736, 0, 4095, 0, 0),
		(drawing, 3737, 0, 4095, 0, 0),
		(drawing, 3738, 0, 4095, 0, 0),
		(drawing, 3739, 0, 4095, 0, 0),
		(drawing, 3740, 0, 4095, 0, 0),
		(drawing, 3741, 0, 4095, 0, 0),
		(drawing, 3742, 0, 4095, 0, 0),
		(drawing, 3743, 0, 4095, 0, 0),
		(drawing, 3744, 0, 4095, 0, 0),
		(drawing, 3745, 0, 4095, 0, 0),
		(drawing, 3746, 0, 4095, 0, 0),
		(drawing, 3747, 0, 4095, 0, 0),
		(drawing, 3748, 0, 4095, 0, 0),
		(drawing, 3749, 0, 4095, 0, 0),
		(drawing, 3750, 0, 4095, 0, 0),
		(drawing, 3751, 0, 4095, 0, 0),
		(drawing, 3752, 0, 4095, 0, 0),
		(drawing, 3753, 0, 4095, 0, 0),
		(drawing, 3754, 0, 4095, 0, 0),
		(drawing, 3755, 0, 4095, 0, 0),
		(drawing, 3756, 0, 4095, 0, 0),
		(drawing, 3757, 0, 4095, 0, 0),
		(drawing, 3758, 0, 4095, 0, 0),
		(drawing, 3759, 0, 4095, 0, 0),
		(drawing, 3760, 0, 4095, 0, 0),
		(drawing, 3761, 0, 4095, 0, 0),
		(drawing, 3762, 0, 4095, 0, 0),
		(drawing, 3763, 0, 4095, 0, 0),
		(drawing, 3764, 0, 4095, 0, 0),
		(drawing, 3765, 0, 4095, 0, 0),
		(drawing, 3766, 0, 4095, 0, 0),
		(drawing, 3767, 0, 4095, 0, 0),
		(drawing, 3768, 0, 4095, 0, 0),
		(drawing, 3769, 0, 4095, 0, 0),
		(drawing, 3770, 0, 4095, 0, 0),
		(drawing, 3771, 0, 4095, 0, 0),
		(drawing, 3772, 0, 4095, 0, 0),
		(drawing, 3773, 0, 4095, 0, 0),
		(drawing, 3774, 0, 4095, 0, 0),
		(drawing, 3775, 0, 4095, 0, 0),
		(drawing, 3776, 0, 4095, 0, 0),
		(drawing, 3777, 0, 4095, 0, 0),
		(drawing, 3778, 0, 4095, 0, 0),
		(drawing, 3779, 0, 4095, 0, 0),
		(drawing, 3780, 0, 4095, 0, 0),
		(drawing, 3781, 0, 4095, 0, 0),
		(drawing, 3782, 0, 4095, 0, 0),
		(drawing, 3783, 0, 4095, 0, 0),
		(drawing, 3784, 0, 4095, 0, 0),
		(drawing, 3785, 0, 4095, 0, 0),
		(drawing, 3786, 0, 4095, 0, 0),
		(drawing, 3787, 0, 4095, 0, 0),
		(drawing, 3788, 0, 4095, 0, 0),
		(drawing, 3789, 0, 4095, 0, 0),
		(drawing, 3790, 0, 4095, 0, 0),
		(drawing, 3791, 0, 4095, 0, 0),
		(drawing, 3792, 0, 4095, 0, 0),
		(drawing, 3793, 0, 4095, 0, 0),
		(drawing, 3794, 0, 4095, 0, 0),
		(drawing, 3795, 0, 4095, 0, 0),
		(drawing, 3796, 0, 4095, 0, 0),
		(drawing, 3797, 0, 4095, 0, 0),
		(drawing, 3798, 0, 4095, 0, 0),
		(drawing, 3799, 0, 4095, 0, 0),
		(drawing, 3800, 0, 4095, 0, 0),
		(drawing, 3801, 0, 4095, 0, 0),
		(drawing, 3802, 0, 4095, 0, 0),
		(drawing, 3803, 0, 4095, 0, 0),
		(drawing, 3804, 0, 4095, 0, 0),
		(drawing, 3805, 0, 4095, 0, 0),
		(drawing, 3806, 0, 4095, 0, 0),
		(drawing, 3807, 0, 4095, 0, 0),
		(drawing, 3808, 0, 4095, 0, 0),
		(drawing, 3809, 0, 4095, 0, 0),
		(drawing, 3810, 0, 4095, 0, 0),
		(drawing, 3811, 0, 4095, 0, 0),
		(drawing, 3812, 0, 4095, 0, 0),
		(drawing, 3813, 0, 4095, 0, 0),
		(drawing, 3814, 0, 4095, 0, 0),
		(drawing, 3815, 0, 4095, 0, 0),
		(drawing, 3816, 0, 4095, 0, 0),
		(drawing, 3817, 0, 4095, 0, 0),
		(drawing, 3818, 0, 4095, 0, 0),
		(drawing, 3819, 0, 4095, 0, 0),
		(drawing, 3820, 0, 4095, 0, 0),
		(drawing, 3821, 0, 4095, 0, 0),
		(drawing, 3822, 0, 4095, 0, 0),
		(drawing, 3823, 0, 4095, 0, 0),
		(drawing, 3824, 0, 4095, 0, 0),
		(drawing, 3825, 0, 4095, 0, 0),
		(drawing, 3826, 0, 4095, 0, 0),
		(drawing, 3827, 0, 4095, 0, 0),
		(drawing, 3828, 0, 4095, 0, 0),
		(drawing, 3829, 0, 4095, 0, 0),
		(drawing, 3830, 0, 4095, 0, 0),
		(drawing, 3831, 0, 4095, 0, 0),
		(drawing, 3832, 0, 4095, 0, 0),
		(drawing, 3833, 0, 4095, 0, 0),
		(drawing, 3834, 0, 4095, 0, 0),
		(drawing, 3835, 0, 4095, 0, 0),
		(drawing, 3836, 0, 4095, 0, 0),
		(drawing, 3837, 0, 4095, 0, 0),
		(drawing, 3838, 0, 4095, 0, 0),
		(drawing, 3839, 0, 4095, 0, 0),
		(drawing, 3840, 0, 4095, 0, 0),
		(drawing, 3841, 0, 4095, 0, 0),
		(drawing, 3842, 0, 4095, 0, 0),
		(drawing, 3843, 0, 4095, 0, 0),
		(drawing, 3844, 0, 4095, 0, 0),
		(drawing, 3845, 0, 4095, 0, 0),
		(drawing, 3846, 0, 4095, 0, 0),
		(drawing, 3847, 0, 4095, 0, 0),
		(drawing, 3848, 0, 4095, 0, 0),
		(drawing, 3849, 0, 4095, 0, 0),
		(drawing, 3850, 0, 4095, 0, 0),
		(drawing, 3851, 0, 4095, 0, 0),
		(drawing, 3852, 0, 4095, 0, 0),
		(drawing, 3853, 0, 4095, 0, 0),
		(drawing, 3854, 0, 4095, 0, 0),
		(drawing, 3855, 0, 4095, 0, 0),
		(drawing, 3856, 0, 4095, 0, 0),
		(drawing, 3857, 0, 4095, 0, 0),
		(drawing, 3858, 0, 4095, 0, 0),
		(drawing, 3859, 0, 4095, 0, 0),
		(drawing, 3860, 0, 4095, 0, 0),
		(drawing, 3861, 0, 4095, 0, 0),
		(drawing, 3862, 0, 4095, 0, 0),
		(drawing, 3863, 0, 4095, 0, 0),
		(drawing, 3864, 0, 4095, 0, 0),
		(drawing, 3865, 0, 4095, 0, 0),
		(drawing, 3866, 0, 4095, 0, 0),
		(drawing, 3867, 0, 4095, 0, 0),
		(drawing, 3868, 0, 4095, 0, 0),
		(drawing, 3869, 0, 4095, 0, 0),
		(drawing, 3870, 0, 4095, 0, 0),
		(drawing, 3871, 0, 4095, 0, 0),
		(drawing, 3872, 0, 4095, 0, 0),
		(drawing, 3873, 0, 4095, 0, 0),
		(drawing, 3874, 0, 4095, 0, 0),
		(drawing, 3875, 0, 4095, 0, 0),
		(drawing, 3876, 0, 4095, 0, 0),
		(drawing, 3877, 0, 4095, 0, 0),
		(drawing, 3878, 0, 4095, 0, 0),
		(drawing, 3879, 0, 4095, 0, 0),
		(drawing, 3880, 0, 4095, 0, 0),
		(drawing, 3881, 0, 4095, 0, 0),
		(drawing, 3882, 0, 4095, 0, 0),
		(drawing, 3883, 0, 4095, 0, 0),
		(drawing, 3884, 0, 4095, 0, 0),
		(drawing, 3885, 0, 4095, 0, 0),
		(drawing, 3886, 0, 4095, 0, 0),
		(drawing, 3887, 0, 4095, 0, 0),
		(drawing, 3888, 0, 4095, 0, 0),
		(drawing, 3889, 0, 4095, 0, 0),
		(drawing, 3890, 0, 4095, 0, 0),
		(drawing, 3891, 0, 4095, 0, 0),
		(drawing, 3892, 0, 4095, 0, 0),
		(drawing, 3893, 0, 4095, 0, 0),
		(drawing, 3894, 0, 4095, 0, 0),
		(drawing, 3895, 0, 4095, 0, 0),
		(drawing, 3896, 0, 4095, 0, 0),
		(drawing, 3897, 0, 4095, 0, 0),
		(drawing, 3898, 0, 4095, 0, 0),
		(drawing, 3899, 0, 4095, 0, 0),
		(drawing, 3900, 0, 4095, 0, 0),
		(drawing, 3901, 0, 4095, 0, 0),
		(drawing, 3902, 0, 4095, 0, 0),
		(drawing, 3903, 0, 4095, 0, 0),
		(drawing, 3904, 0, 4095, 0, 0),
		(drawing, 3905, 0, 4095, 0, 0),
		(drawing, 3906, 0, 4095, 0, 0),
		(drawing, 3907, 0, 4095, 0, 0),
		(drawing, 3908, 0, 4095, 0, 0),
		(drawing, 3909, 0, 4095, 0, 0),
		(drawing, 3910, 0, 4095, 0, 0),
		(drawing, 3911, 0, 4095, 0, 0),
		(drawing, 3912, 0, 4095, 0, 0),
		(drawing, 3913, 0, 4095, 0, 0),
		(drawing, 3914, 0, 4095, 0, 0),
		(drawing, 3915, 0, 4095, 0, 0),
		(drawing, 3916, 0, 4095, 0, 0),
		(drawing, 3917, 0, 4095, 0, 0),
		(drawing, 3918, 0, 4095, 0, 0),
		(drawing, 3919, 0, 4095, 0, 0),
		(drawing, 3920, 0, 4095, 0, 0),
		(drawing, 3921, 0, 4095, 0, 0),
		(drawing, 3922, 0, 4095, 0, 0),
		(drawing, 3923, 0, 4095, 0, 0),
		(drawing, 3924, 0, 4095, 0, 0),
		(drawing, 3925, 0, 4095, 0, 0),
		(drawing, 3926, 0, 4095, 0, 0),
		(drawing, 3927, 0, 4095, 0, 0),
		(drawing, 3928, 0, 4095, 0, 0),
		(drawing, 3929, 0, 4095, 0, 0),
		(drawing, 3930, 0, 4095, 0, 0),
		(drawing, 3931, 0, 4095, 0, 0),
		(drawing, 3932, 0, 4095, 0, 0),
		(drawing, 3933, 0, 4095, 0, 0),
		(drawing, 3934, 0, 4095, 0, 0),
		(drawing, 3935, 0, 4095, 0, 0),
		(drawing, 3936, 0, 4095, 0, 0),
		(drawing, 3937, 0, 4095, 0, 0),
		(drawing, 3938, 0, 4095, 0, 0),
		(drawing, 3939, 0, 4095, 0, 0),
		(drawing, 3940, 0, 4095, 0, 0),
		(drawing, 3941, 0, 4095, 0, 0),
		(drawing, 3942, 0, 4095, 0, 0),
		(drawing, 3943, 0, 4095, 0, 0),
		(drawing, 3944, 0, 4095, 0, 0),
		(drawing, 3945, 0, 4095, 0, 0),
		(drawing, 3946, 0, 4095, 0, 0),
		(drawing, 3947, 0, 4095, 0, 0),
		(drawing, 3948, 0, 4095, 0, 0),
		(drawing, 3949, 0, 4095, 0, 0),
		(drawing, 3950, 0, 4095, 0, 0),
		(drawing, 3951, 0, 4095, 0, 0),
		(drawing, 3952, 0, 4095, 0, 0),
		(drawing, 3953, 0, 4095, 0, 0),
		(drawing, 3954, 0, 4095, 0, 0),
		(drawing, 3955, 0, 4095, 0, 0),
		(drawing, 3956, 0, 4095, 0, 0),
		(drawing, 3957, 0, 4095, 0, 0),
		(drawing, 3958, 0, 4095, 0, 0),
		(drawing, 3959, 0, 4095, 0, 0),
		(drawing, 3960, 0, 4095, 0, 0),
		(drawing, 3961, 0, 4095, 0, 0),
		(drawing, 3962, 0, 4095, 0, 0),
		(drawing, 3963, 0, 4095, 0, 0),
		(drawing, 3964, 0, 4095, 0, 0),
		(drawing, 3965, 0, 4095, 0, 0),
		(drawing, 3966, 0, 4095, 0, 0),
		(drawing, 3967, 0, 4095, 0, 0),
		(drawing, 3968, 0, 4095, 0, 0),
		(drawing, 3969, 0, 4095, 0, 0),
		(drawing, 3970, 0, 4095, 0, 0),
		(drawing, 3971, 0, 4095, 0, 0),
		(drawing, 3972, 0, 4095, 0, 0),
		(drawing, 3973, 0, 4095, 0, 0),
		(drawing, 3974, 0, 4095, 0, 0),
		(drawing, 3975, 0, 4095, 0, 0),
		(drawing, 3976, 0, 4095, 0, 0),
		(drawing, 3977, 0, 4095, 0, 0),
		(drawing, 3978, 0, 4095, 0, 0),
		(drawing, 3979, 0, 4095, 0, 0),
		(drawing, 3980, 0, 4095, 0, 0),
		(drawing, 3981, 0, 4095, 0, 0),
		(drawing, 3982, 0, 4095, 0, 0),
		(drawing, 3983, 0, 4095, 0, 0),
		(drawing, 3984, 0, 4095, 0, 0),
		(drawing, 3985, 0, 4095, 0, 0),
		(drawing, 3986, 0, 4095, 0, 0),
		(drawing, 3987, 0, 4095, 0, 0),
		(drawing, 3988, 0, 4095, 0, 0),
		(drawing, 3989, 0, 4095, 0, 0),
		(drawing, 3990, 0, 4095, 0, 0),
		(drawing, 3991, 0, 4095, 0, 0),
		(drawing, 3992, 0, 4095, 0, 0),
		(drawing, 3993, 0, 4095, 0, 0),
		(drawing, 3994, 0, 4095, 0, 0),
		(drawing, 3995, 0, 4095, 0, 0),
		(drawing, 3996, 0, 4095, 0, 0),
		(drawing, 3997, 0, 4095, 0, 0),
		(drawing, 3998, 0, 4095, 0, 0),
		(drawing, 3999, 0, 4095, 0, 0),
		(drawing, 4000, 0, 4095, 0, 0),
		(drawing, 4001, 0, 4095, 0, 0),
		(drawing, 4002, 0, 4095, 0, 0),
		(drawing, 4003, 0, 4095, 0, 0),
		(drawing, 4004, 0, 4095, 0, 0),
		(drawing, 4005, 0, 4095, 0, 0),
		(drawing, 4006, 0, 4095, 0, 0),
		(drawing, 4007, 0, 4095, 0, 0),
		(drawing, 4008, 0, 4095, 0, 0),
		(drawing, 4009, 0, 4095, 0, 0),
		(drawing, 4010, 0, 4095, 0, 0),
		(drawing, 4011, 0, 4095, 0, 0),
		(drawing, 4012, 0, 4095, 0, 0),
		(drawing, 4013, 0, 4095, 0, 0),
		(drawing, 4014, 0, 4095, 0, 0),
		(drawing, 4015, 0, 4095, 0, 0),
		(drawing, 4016, 0, 4095, 0, 0),
		(drawing, 4017, 0, 4095, 0, 0),
		(drawing, 4018, 0, 4095, 0, 0),
		(drawing, 4019, 0, 4095, 0, 0),
		(drawing, 4020, 0, 4095, 0, 0),
		(drawing, 4021, 0, 4095, 0, 0),
		(drawing, 4022, 0, 4095, 0, 0),
		(drawing, 4023, 0, 4095, 0, 0),
		(drawing, 4024, 0, 4095, 0, 0),
		(drawing, 4025, 0, 4095, 0, 0),
		(drawing, 4026, 0, 4095, 0, 0),
		(drawing, 4027, 0, 4095, 0, 0),
		(drawing, 4028, 0, 4095, 0, 0),
		(drawing, 4029, 0, 4095, 0, 0),
		(drawing, 4030, 0, 4095, 0, 0),
		(drawing, 4031, 0, 4095, 0, 0),
		(drawing, 4032, 0, 4095, 0, 0),
		(drawing, 4033, 0, 4095, 0, 0),
		(drawing, 4034, 0, 4095, 0, 0),
		(drawing, 4035, 0, 4095, 0, 0),
		(drawing, 4036, 0, 4095, 0, 0),
		(drawing, 4037, 0, 4095, 0, 0),
		(drawing, 4038, 0, 4095, 0, 0),
		(drawing, 4039, 0, 4095, 0, 0),
		(drawing, 4040, 0, 4095, 0, 0),
		(drawing, 4041, 0, 4095, 0, 0),
		(drawing, 4042, 0, 4095, 0, 0),
		(drawing, 4043, 0, 4095, 0, 0),
		(drawing, 4044, 0, 4095, 0, 0),
		(drawing, 4045, 0, 4095, 0, 0),
		(drawing, 4046, 0, 4095, 0, 0),
		(drawing, 4047, 0, 4095, 0, 0),
		(drawing, 4048, 0, 4095, 0, 0),
		(drawing, 4049, 0, 4095, 0, 0),
		(drawing, 4050, 0, 4095, 0, 0),
		(drawing, 4051, 0, 4095, 0, 0),
		(drawing, 4052, 0, 4095, 0, 0),
		(drawing, 4053, 0, 4095, 0, 0),
		(drawing, 4054, 0, 4095, 0, 0),
		(drawing, 4055, 0, 4095, 0, 0),
		(drawing, 4056, 0, 4095, 0, 0),
		(drawing, 4057, 0, 4095, 0, 0),
		(drawing, 4058, 0, 4095, 0, 0),
		(drawing, 4059, 0, 4095, 0, 0),
		(drawing, 4060, 0, 4095, 0, 0),
		(drawing, 4061, 0, 4095, 0, 0),
		(drawing, 4062, 0, 4095, 0, 0),
		(drawing, 4063, 0, 4095, 0, 0),
		(drawing, 4064, 0, 4095, 0, 0),
		(drawing, 4065, 0, 4095, 0, 0),
		(drawing, 4066, 0, 4095, 0, 0),
		(drawing, 4067, 0, 4095, 0, 0),
		(drawing, 4068, 0, 4095, 0, 0),
		(drawing, 4069, 0, 4095, 0, 0),
		(drawing, 4070, 0, 4095, 0, 0),
		(drawing, 4071, 0, 4095, 0, 0),
		(drawing, 4072, 0, 4095, 0, 0),
		(drawing, 4073, 0, 4095, 0, 0),
		(drawing, 4074, 0, 4095, 0, 0),
		(drawing, 4075, 0, 4095, 0, 0),
		(drawing, 4076, 0, 4095, 0, 0),
		(drawing, 4077, 0, 4095, 0, 0),
		(drawing, 4078, 0, 4095, 0, 0),
		(drawing, 4079, 0, 4095, 0, 0),
		(drawing, 4080, 0, 4095, 0, 0),
		(drawing, 4081, 0, 4095, 0, 0),
		(drawing, 4082, 0, 4095, 0, 0),
		(drawing, 4083, 0, 4095, 0, 0),
		(drawing, 4084, 0, 4095, 0, 0),
		(drawing, 4085, 0, 4095, 0, 0),
		(drawing, 4086, 0, 4095, 0, 0),
		(drawing, 4087, 0, 4095, 0, 0),
		(drawing, 4088, 0, 4095, 0, 0),
		(drawing, 4089, 0, 4095, 0, 0),
		(drawing, 4090, 0, 4095, 0, 0),
		(drawing, 4091, 0, 4095, 0, 0),
		(drawing, 4092, 0, 4095, 0, 0),
		(drawing, 4093, 0, 4095, 0, 0),
		(drawing, 4094, 0, 4095, 0, 0),
		(done, 4095, 0, 4095, 0, 0)
	);
END PACKAGE ex1_data_pak;
