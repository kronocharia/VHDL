-- advanced test 7
-- draw line from (0,0) to (2048,30)
-- testing the calculation of err1 and err2 with large number (number larger or equal to 2048) 
-- and also the comparison of err1 and err2.

PACKAGE ex1_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 0, 0, 0),
		(start, 0, 0, 2048, 30, 0),
		(drawing, 0, 0, 2048, 30, 0),
		(drawing, 1, 0, 2048, 30, 0),
		(drawing, 2, 0, 2048, 30, 0),
		(drawing, 3, 0, 2048, 30, 0),
		(drawing, 4, 0, 2048, 30, 0),
		(drawing, 5, 0, 2048, 30, 0),
		(drawing, 6, 0, 2048, 30, 0),
		(drawing, 7, 0, 2048, 30, 0),
		(drawing, 8, 0, 2048, 30, 0),
		(drawing, 9, 0, 2048, 30, 0),
		(drawing, 10, 0, 2048, 30, 0),
		(drawing, 11, 0, 2048, 30, 0),
		(drawing, 12, 0, 2048, 30, 0),
		(drawing, 13, 0, 2048, 30, 0),
		(drawing, 14, 0, 2048, 30, 0),
		(drawing, 15, 0, 2048, 30, 0),
		(drawing, 16, 0, 2048, 30, 0),
		(drawing, 17, 0, 2048, 30, 0),
		(drawing, 18, 0, 2048, 30, 0),
		(drawing, 19, 0, 2048, 30, 0),
		(drawing, 20, 0, 2048, 30, 0),
		(drawing, 21, 0, 2048, 30, 0),
		(drawing, 22, 0, 2048, 30, 0),
		(drawing, 23, 0, 2048, 30, 0),
		(drawing, 24, 0, 2048, 30, 0),
		(drawing, 25, 0, 2048, 30, 0),
		(drawing, 26, 0, 2048, 30, 0),
		(drawing, 27, 0, 2048, 30, 0),
		(drawing, 28, 0, 2048, 30, 0),
		(drawing, 29, 0, 2048, 30, 0),
		(drawing, 30, 0, 2048, 30, 0),
		(drawing, 31, 0, 2048, 30, 0),
		(drawing, 32, 0, 2048, 30, 0),
		(drawing, 33, 0, 2048, 30, 0),
		(drawing, 34, 0, 2048, 30, 0),
		(drawing, 35, 1, 2048, 30, 0),
		(drawing, 36, 1, 2048, 30, 0),
		(drawing, 37, 1, 2048, 30, 0),
		(drawing, 38, 1, 2048, 30, 0),
		(drawing, 39, 1, 2048, 30, 0),
		(drawing, 40, 1, 2048, 30, 0),
		(drawing, 41, 1, 2048, 30, 0),
		(drawing, 42, 1, 2048, 30, 0),
		(drawing, 43, 1, 2048, 30, 0),
		(drawing, 44, 1, 2048, 30, 0),
		(drawing, 45, 1, 2048, 30, 0),
		(drawing, 46, 1, 2048, 30, 0),
		(drawing, 47, 1, 2048, 30, 0),
		(drawing, 48, 1, 2048, 30, 0),
		(drawing, 49, 1, 2048, 30, 0),
		(drawing, 50, 1, 2048, 30, 0),
		(drawing, 51, 1, 2048, 30, 0),
		(drawing, 52, 1, 2048, 30, 0),
		(drawing, 53, 1, 2048, 30, 0),
		(drawing, 54, 1, 2048, 30, 0),
		(drawing, 55, 1, 2048, 30, 0),
		(drawing, 56, 1, 2048, 30, 0),
		(drawing, 57, 1, 2048, 30, 0),
		(drawing, 58, 1, 2048, 30, 0),
		(drawing, 59, 1, 2048, 30, 0),
		(drawing, 60, 1, 2048, 30, 0),
		(drawing, 61, 1, 2048, 30, 0),
		(drawing, 62, 1, 2048, 30, 0),
		(drawing, 63, 1, 2048, 30, 0),
		(drawing, 64, 1, 2048, 30, 0),
		(drawing, 65, 1, 2048, 30, 0),
		(drawing, 66, 1, 2048, 30, 0),
		(drawing, 67, 1, 2048, 30, 0),
		(drawing, 68, 1, 2048, 30, 0),
		(drawing, 69, 1, 2048, 30, 0),
		(drawing, 70, 1, 2048, 30, 0),
		(drawing, 71, 1, 2048, 30, 0),
		(drawing, 72, 1, 2048, 30, 0),
		(drawing, 73, 1, 2048, 30, 0),
		(drawing, 74, 1, 2048, 30, 0),
		(drawing, 75, 1, 2048, 30, 0),
		(drawing, 76, 1, 2048, 30, 0),
		(drawing, 77, 1, 2048, 30, 0),
		(drawing, 78, 1, 2048, 30, 0),
		(drawing, 79, 1, 2048, 30, 0),
		(drawing, 80, 1, 2048, 30, 0),
		(drawing, 81, 1, 2048, 30, 0),
		(drawing, 82, 1, 2048, 30, 0),
		(drawing, 83, 1, 2048, 30, 0),
		(drawing, 84, 1, 2048, 30, 0),
		(drawing, 85, 1, 2048, 30, 0),
		(drawing, 86, 1, 2048, 30, 0),
		(drawing, 87, 1, 2048, 30, 0),
		(drawing, 88, 1, 2048, 30, 0),
		(drawing, 89, 1, 2048, 30, 0),
		(drawing, 90, 1, 2048, 30, 0),
		(drawing, 91, 1, 2048, 30, 0),
		(drawing, 92, 1, 2048, 30, 0),
		(drawing, 93, 1, 2048, 30, 0),
		(drawing, 94, 1, 2048, 30, 0),
		(drawing, 95, 1, 2048, 30, 0),
		(drawing, 96, 1, 2048, 30, 0),
		(drawing, 97, 1, 2048, 30, 0),
		(drawing, 98, 1, 2048, 30, 0),
		(drawing, 99, 1, 2048, 30, 0),
		(drawing, 100, 1, 2048, 30, 0),
		(drawing, 101, 1, 2048, 30, 0),
		(drawing, 102, 1, 2048, 30, 0),
		(drawing, 103, 2, 2048, 30, 0),
		(drawing, 104, 2, 2048, 30, 0),
		(drawing, 105, 2, 2048, 30, 0),
		(drawing, 106, 2, 2048, 30, 0),
		(drawing, 107, 2, 2048, 30, 0),
		(drawing, 108, 2, 2048, 30, 0),
		(drawing, 109, 2, 2048, 30, 0),
		(drawing, 110, 2, 2048, 30, 0),
		(drawing, 111, 2, 2048, 30, 0),
		(drawing, 112, 2, 2048, 30, 0),
		(drawing, 113, 2, 2048, 30, 0),
		(drawing, 114, 2, 2048, 30, 0),
		(drawing, 115, 2, 2048, 30, 0),
		(drawing, 116, 2, 2048, 30, 0),
		(drawing, 117, 2, 2048, 30, 0),
		(drawing, 118, 2, 2048, 30, 0),
		(drawing, 119, 2, 2048, 30, 0),
		(drawing, 120, 2, 2048, 30, 0),
		(drawing, 121, 2, 2048, 30, 0),
		(drawing, 122, 2, 2048, 30, 0),
		(drawing, 123, 2, 2048, 30, 0),
		(drawing, 124, 2, 2048, 30, 0),
		(drawing, 125, 2, 2048, 30, 0),
		(drawing, 126, 2, 2048, 30, 0),
		(drawing, 127, 2, 2048, 30, 0),
		(drawing, 128, 2, 2048, 30, 0),
		(drawing, 129, 2, 2048, 30, 0),
		(drawing, 130, 2, 2048, 30, 0),
		(drawing, 131, 2, 2048, 30, 0),
		(drawing, 132, 2, 2048, 30, 0),
		(drawing, 133, 2, 2048, 30, 0),
		(drawing, 134, 2, 2048, 30, 0),
		(drawing, 135, 2, 2048, 30, 0),
		(drawing, 136, 2, 2048, 30, 0),
		(drawing, 137, 2, 2048, 30, 0),
		(drawing, 138, 2, 2048, 30, 0),
		(drawing, 139, 2, 2048, 30, 0),
		(drawing, 140, 2, 2048, 30, 0),
		(drawing, 141, 2, 2048, 30, 0),
		(drawing, 142, 2, 2048, 30, 0),
		(drawing, 143, 2, 2048, 30, 0),
		(drawing, 144, 2, 2048, 30, 0),
		(drawing, 145, 2, 2048, 30, 0),
		(drawing, 146, 2, 2048, 30, 0),
		(drawing, 147, 2, 2048, 30, 0),
		(drawing, 148, 2, 2048, 30, 0),
		(drawing, 149, 2, 2048, 30, 0),
		(drawing, 150, 2, 2048, 30, 0),
		(drawing, 151, 2, 2048, 30, 0),
		(drawing, 152, 2, 2048, 30, 0),
		(drawing, 153, 2, 2048, 30, 0),
		(drawing, 154, 2, 2048, 30, 0),
		(drawing, 155, 2, 2048, 30, 0),
		(drawing, 156, 2, 2048, 30, 0),
		(drawing, 157, 2, 2048, 30, 0),
		(drawing, 158, 2, 2048, 30, 0),
		(drawing, 159, 2, 2048, 30, 0),
		(drawing, 160, 2, 2048, 30, 0),
		(drawing, 161, 2, 2048, 30, 0),
		(drawing, 162, 2, 2048, 30, 0),
		(drawing, 163, 2, 2048, 30, 0),
		(drawing, 164, 2, 2048, 30, 0),
		(drawing, 165, 2, 2048, 30, 0),
		(drawing, 166, 2, 2048, 30, 0),
		(drawing, 167, 2, 2048, 30, 0),
		(drawing, 168, 2, 2048, 30, 0),
		(drawing, 169, 2, 2048, 30, 0),
		(drawing, 170, 2, 2048, 30, 0),
		(drawing, 171, 3, 2048, 30, 0),
		(drawing, 172, 3, 2048, 30, 0),
		(drawing, 173, 3, 2048, 30, 0),
		(drawing, 174, 3, 2048, 30, 0),
		(drawing, 175, 3, 2048, 30, 0),
		(drawing, 176, 3, 2048, 30, 0),
		(drawing, 177, 3, 2048, 30, 0),
		(drawing, 178, 3, 2048, 30, 0),
		(drawing, 179, 3, 2048, 30, 0),
		(drawing, 180, 3, 2048, 30, 0),
		(drawing, 181, 3, 2048, 30, 0),
		(drawing, 182, 3, 2048, 30, 0),
		(drawing, 183, 3, 2048, 30, 0),
		(drawing, 184, 3, 2048, 30, 0),
		(drawing, 185, 3, 2048, 30, 0),
		(drawing, 186, 3, 2048, 30, 0),
		(drawing, 187, 3, 2048, 30, 0),
		(drawing, 188, 3, 2048, 30, 0),
		(drawing, 189, 3, 2048, 30, 0),
		(drawing, 190, 3, 2048, 30, 0),
		(drawing, 191, 3, 2048, 30, 0),
		(drawing, 192, 3, 2048, 30, 0),
		(drawing, 193, 3, 2048, 30, 0),
		(drawing, 194, 3, 2048, 30, 0),
		(drawing, 195, 3, 2048, 30, 0),
		(drawing, 196, 3, 2048, 30, 0),
		(drawing, 197, 3, 2048, 30, 0),
		(drawing, 198, 3, 2048, 30, 0),
		(drawing, 199, 3, 2048, 30, 0),
		(drawing, 200, 3, 2048, 30, 0),
		(drawing, 201, 3, 2048, 30, 0),
		(drawing, 202, 3, 2048, 30, 0),
		(drawing, 203, 3, 2048, 30, 0),
		(drawing, 204, 3, 2048, 30, 0),
		(drawing, 205, 3, 2048, 30, 0),
		(drawing, 206, 3, 2048, 30, 0),
		(drawing, 207, 3, 2048, 30, 0),
		(drawing, 208, 3, 2048, 30, 0),
		(drawing, 209, 3, 2048, 30, 0),
		(drawing, 210, 3, 2048, 30, 0),
		(drawing, 211, 3, 2048, 30, 0),
		(drawing, 212, 3, 2048, 30, 0),
		(drawing, 213, 3, 2048, 30, 0),
		(drawing, 214, 3, 2048, 30, 0),
		(drawing, 215, 3, 2048, 30, 0),
		(drawing, 216, 3, 2048, 30, 0),
		(drawing, 217, 3, 2048, 30, 0),
		(drawing, 218, 3, 2048, 30, 0),
		(drawing, 219, 3, 2048, 30, 0),
		(drawing, 220, 3, 2048, 30, 0),
		(drawing, 221, 3, 2048, 30, 0),
		(drawing, 222, 3, 2048, 30, 0),
		(drawing, 223, 3, 2048, 30, 0),
		(drawing, 224, 3, 2048, 30, 0),
		(drawing, 225, 3, 2048, 30, 0),
		(drawing, 226, 3, 2048, 30, 0),
		(drawing, 227, 3, 2048, 30, 0),
		(drawing, 228, 3, 2048, 30, 0),
		(drawing, 229, 3, 2048, 30, 0),
		(drawing, 230, 3, 2048, 30, 0),
		(drawing, 231, 3, 2048, 30, 0),
		(drawing, 232, 3, 2048, 30, 0),
		(drawing, 233, 3, 2048, 30, 0),
		(drawing, 234, 3, 2048, 30, 0),
		(drawing, 235, 3, 2048, 30, 0),
		(drawing, 236, 3, 2048, 30, 0),
		(drawing, 237, 3, 2048, 30, 0),
		(drawing, 238, 3, 2048, 30, 0),
		(drawing, 239, 4, 2048, 30, 0),
		(drawing, 240, 4, 2048, 30, 0),
		(drawing, 241, 4, 2048, 30, 0),
		(drawing, 242, 4, 2048, 30, 0),
		(drawing, 243, 4, 2048, 30, 0),
		(drawing, 244, 4, 2048, 30, 0),
		(drawing, 245, 4, 2048, 30, 0),
		(drawing, 246, 4, 2048, 30, 0),
		(drawing, 247, 4, 2048, 30, 0),
		(drawing, 248, 4, 2048, 30, 0),
		(drawing, 249, 4, 2048, 30, 0),
		(drawing, 250, 4, 2048, 30, 0),
		(drawing, 251, 4, 2048, 30, 0),
		(drawing, 252, 4, 2048, 30, 0),
		(drawing, 253, 4, 2048, 30, 0),
		(drawing, 254, 4, 2048, 30, 0),
		(drawing, 255, 4, 2048, 30, 0),
		(drawing, 256, 4, 2048, 30, 0),
		(drawing, 257, 4, 2048, 30, 0),
		(drawing, 258, 4, 2048, 30, 0),
		(drawing, 259, 4, 2048, 30, 0),
		(drawing, 260, 4, 2048, 30, 0),
		(drawing, 261, 4, 2048, 30, 0),
		(drawing, 262, 4, 2048, 30, 0),
		(drawing, 263, 4, 2048, 30, 0),
		(drawing, 264, 4, 2048, 30, 0),
		(drawing, 265, 4, 2048, 30, 0),
		(drawing, 266, 4, 2048, 30, 0),
		(drawing, 267, 4, 2048, 30, 0),
		(drawing, 268, 4, 2048, 30, 0),
		(drawing, 269, 4, 2048, 30, 0),
		(drawing, 270, 4, 2048, 30, 0),
		(drawing, 271, 4, 2048, 30, 0),
		(drawing, 272, 4, 2048, 30, 0),
		(drawing, 273, 4, 2048, 30, 0),
		(drawing, 274, 4, 2048, 30, 0),
		(drawing, 275, 4, 2048, 30, 0),
		(drawing, 276, 4, 2048, 30, 0),
		(drawing, 277, 4, 2048, 30, 0),
		(drawing, 278, 4, 2048, 30, 0),
		(drawing, 279, 4, 2048, 30, 0),
		(drawing, 280, 4, 2048, 30, 0),
		(drawing, 281, 4, 2048, 30, 0),
		(drawing, 282, 4, 2048, 30, 0),
		(drawing, 283, 4, 2048, 30, 0),
		(drawing, 284, 4, 2048, 30, 0),
		(drawing, 285, 4, 2048, 30, 0),
		(drawing, 286, 4, 2048, 30, 0),
		(drawing, 287, 4, 2048, 30, 0),
		(drawing, 288, 4, 2048, 30, 0),
		(drawing, 289, 4, 2048, 30, 0),
		(drawing, 290, 4, 2048, 30, 0),
		(drawing, 291, 4, 2048, 30, 0),
		(drawing, 292, 4, 2048, 30, 0),
		(drawing, 293, 4, 2048, 30, 0),
		(drawing, 294, 4, 2048, 30, 0),
		(drawing, 295, 4, 2048, 30, 0),
		(drawing, 296, 4, 2048, 30, 0),
		(drawing, 297, 4, 2048, 30, 0),
		(drawing, 298, 4, 2048, 30, 0),
		(drawing, 299, 4, 2048, 30, 0),
		(drawing, 300, 4, 2048, 30, 0),
		(drawing, 301, 4, 2048, 30, 0),
		(drawing, 302, 4, 2048, 30, 0),
		(drawing, 303, 4, 2048, 30, 0),
		(drawing, 304, 4, 2048, 30, 0),
		(drawing, 305, 4, 2048, 30, 0),
		(drawing, 306, 4, 2048, 30, 0),
		(drawing, 307, 4, 2048, 30, 0),
		(drawing, 308, 5, 2048, 30, 0),
		(drawing, 309, 5, 2048, 30, 0),
		(drawing, 310, 5, 2048, 30, 0),
		(drawing, 311, 5, 2048, 30, 0),
		(drawing, 312, 5, 2048, 30, 0),
		(drawing, 313, 5, 2048, 30, 0),
		(drawing, 314, 5, 2048, 30, 0),
		(drawing, 315, 5, 2048, 30, 0),
		(drawing, 316, 5, 2048, 30, 0),
		(drawing, 317, 5, 2048, 30, 0),
		(drawing, 318, 5, 2048, 30, 0),
		(drawing, 319, 5, 2048, 30, 0),
		(drawing, 320, 5, 2048, 30, 0),
		(drawing, 321, 5, 2048, 30, 0),
		(drawing, 322, 5, 2048, 30, 0),
		(drawing, 323, 5, 2048, 30, 0),
		(drawing, 324, 5, 2048, 30, 0),
		(drawing, 325, 5, 2048, 30, 0),
		(drawing, 326, 5, 2048, 30, 0),
		(drawing, 327, 5, 2048, 30, 0),
		(drawing, 328, 5, 2048, 30, 0),
		(drawing, 329, 5, 2048, 30, 0),
		(drawing, 330, 5, 2048, 30, 0),
		(drawing, 331, 5, 2048, 30, 0),
		(drawing, 332, 5, 2048, 30, 0),
		(drawing, 333, 5, 2048, 30, 0),
		(drawing, 334, 5, 2048, 30, 0),
		(drawing, 335, 5, 2048, 30, 0),
		(drawing, 336, 5, 2048, 30, 0),
		(drawing, 337, 5, 2048, 30, 0),
		(drawing, 338, 5, 2048, 30, 0),
		(drawing, 339, 5, 2048, 30, 0),
		(drawing, 340, 5, 2048, 30, 0),
		(drawing, 341, 5, 2048, 30, 0),
		(drawing, 342, 5, 2048, 30, 0),
		(drawing, 343, 5, 2048, 30, 0),
		(drawing, 344, 5, 2048, 30, 0),
		(drawing, 345, 5, 2048, 30, 0),
		(drawing, 346, 5, 2048, 30, 0),
		(drawing, 347, 5, 2048, 30, 0),
		(drawing, 348, 5, 2048, 30, 0),
		(drawing, 349, 5, 2048, 30, 0),
		(drawing, 350, 5, 2048, 30, 0),
		(drawing, 351, 5, 2048, 30, 0),
		(drawing, 352, 5, 2048, 30, 0),
		(drawing, 353, 5, 2048, 30, 0),
		(drawing, 354, 5, 2048, 30, 0),
		(drawing, 355, 5, 2048, 30, 0),
		(drawing, 356, 5, 2048, 30, 0),
		(drawing, 357, 5, 2048, 30, 0),
		(drawing, 358, 5, 2048, 30, 0),
		(drawing, 359, 5, 2048, 30, 0),
		(drawing, 360, 5, 2048, 30, 0),
		(drawing, 361, 5, 2048, 30, 0),
		(drawing, 362, 5, 2048, 30, 0),
		(drawing, 363, 5, 2048, 30, 0),
		(drawing, 364, 5, 2048, 30, 0),
		(drawing, 365, 5, 2048, 30, 0),
		(drawing, 366, 5, 2048, 30, 0),
		(drawing, 367, 5, 2048, 30, 0),
		(drawing, 368, 5, 2048, 30, 0),
		(drawing, 369, 5, 2048, 30, 0),
		(drawing, 370, 5, 2048, 30, 0),
		(drawing, 371, 5, 2048, 30, 0),
		(drawing, 372, 5, 2048, 30, 0),
		(drawing, 373, 5, 2048, 30, 0),
		(drawing, 374, 5, 2048, 30, 0),
		(drawing, 375, 5, 2048, 30, 0),
		(drawing, 376, 6, 2048, 30, 0),
		(drawing, 377, 6, 2048, 30, 0),
		(drawing, 378, 6, 2048, 30, 0),
		(drawing, 379, 6, 2048, 30, 0),
		(drawing, 380, 6, 2048, 30, 0),
		(drawing, 381, 6, 2048, 30, 0),
		(drawing, 382, 6, 2048, 30, 0),
		(drawing, 383, 6, 2048, 30, 0),
		(drawing, 384, 6, 2048, 30, 0),
		(drawing, 385, 6, 2048, 30, 0),
		(drawing, 386, 6, 2048, 30, 0),
		(drawing, 387, 6, 2048, 30, 0),
		(drawing, 388, 6, 2048, 30, 0),
		(drawing, 389, 6, 2048, 30, 0),
		(drawing, 390, 6, 2048, 30, 0),
		(drawing, 391, 6, 2048, 30, 0),
		(drawing, 392, 6, 2048, 30, 0),
		(drawing, 393, 6, 2048, 30, 0),
		(drawing, 394, 6, 2048, 30, 0),
		(drawing, 395, 6, 2048, 30, 0),
		(drawing, 396, 6, 2048, 30, 0),
		(drawing, 397, 6, 2048, 30, 0),
		(drawing, 398, 6, 2048, 30, 0),
		(drawing, 399, 6, 2048, 30, 0),
		(drawing, 400, 6, 2048, 30, 0),
		(drawing, 401, 6, 2048, 30, 0),
		(drawing, 402, 6, 2048, 30, 0),
		(drawing, 403, 6, 2048, 30, 0),
		(drawing, 404, 6, 2048, 30, 0),
		(drawing, 405, 6, 2048, 30, 0),
		(drawing, 406, 6, 2048, 30, 0),
		(drawing, 407, 6, 2048, 30, 0),
		(drawing, 408, 6, 2048, 30, 0),
		(drawing, 409, 6, 2048, 30, 0),
		(drawing, 410, 6, 2048, 30, 0),
		(drawing, 411, 6, 2048, 30, 0),
		(drawing, 412, 6, 2048, 30, 0),
		(drawing, 413, 6, 2048, 30, 0),
		(drawing, 414, 6, 2048, 30, 0),
		(drawing, 415, 6, 2048, 30, 0),
		(drawing, 416, 6, 2048, 30, 0),
		(drawing, 417, 6, 2048, 30, 0),
		(drawing, 418, 6, 2048, 30, 0),
		(drawing, 419, 6, 2048, 30, 0),
		(drawing, 420, 6, 2048, 30, 0),
		(drawing, 421, 6, 2048, 30, 0),
		(drawing, 422, 6, 2048, 30, 0),
		(drawing, 423, 6, 2048, 30, 0),
		(drawing, 424, 6, 2048, 30, 0),
		(drawing, 425, 6, 2048, 30, 0),
		(drawing, 426, 6, 2048, 30, 0),
		(drawing, 427, 6, 2048, 30, 0),
		(drawing, 428, 6, 2048, 30, 0),
		(drawing, 429, 6, 2048, 30, 0),
		(drawing, 430, 6, 2048, 30, 0),
		(drawing, 431, 6, 2048, 30, 0),
		(drawing, 432, 6, 2048, 30, 0),
		(drawing, 433, 6, 2048, 30, 0),
		(drawing, 434, 6, 2048, 30, 0),
		(drawing, 435, 6, 2048, 30, 0),
		(drawing, 436, 6, 2048, 30, 0),
		(drawing, 437, 6, 2048, 30, 0),
		(drawing, 438, 6, 2048, 30, 0),
		(drawing, 439, 6, 2048, 30, 0),
		(drawing, 440, 6, 2048, 30, 0),
		(drawing, 441, 6, 2048, 30, 0),
		(drawing, 442, 6, 2048, 30, 0),
		(drawing, 443, 6, 2048, 30, 0),
		(drawing, 444, 7, 2048, 30, 0),
		(drawing, 445, 7, 2048, 30, 0),
		(drawing, 446, 7, 2048, 30, 0),
		(drawing, 447, 7, 2048, 30, 0),
		(drawing, 448, 7, 2048, 30, 0),
		(drawing, 449, 7, 2048, 30, 0),
		(drawing, 450, 7, 2048, 30, 0),
		(drawing, 451, 7, 2048, 30, 0),
		(drawing, 452, 7, 2048, 30, 0),
		(drawing, 453, 7, 2048, 30, 0),
		(drawing, 454, 7, 2048, 30, 0),
		(drawing, 455, 7, 2048, 30, 0),
		(drawing, 456, 7, 2048, 30, 0),
		(drawing, 457, 7, 2048, 30, 0),
		(drawing, 458, 7, 2048, 30, 0),
		(drawing, 459, 7, 2048, 30, 0),
		(drawing, 460, 7, 2048, 30, 0),
		(drawing, 461, 7, 2048, 30, 0),
		(drawing, 462, 7, 2048, 30, 0),
		(drawing, 463, 7, 2048, 30, 0),
		(drawing, 464, 7, 2048, 30, 0),
		(drawing, 465, 7, 2048, 30, 0),
		(drawing, 466, 7, 2048, 30, 0),
		(drawing, 467, 7, 2048, 30, 0),
		(drawing, 468, 7, 2048, 30, 0),
		(drawing, 469, 7, 2048, 30, 0),
		(drawing, 470, 7, 2048, 30, 0),
		(drawing, 471, 7, 2048, 30, 0),
		(drawing, 472, 7, 2048, 30, 0),
		(drawing, 473, 7, 2048, 30, 0),
		(drawing, 474, 7, 2048, 30, 0),
		(drawing, 475, 7, 2048, 30, 0),
		(drawing, 476, 7, 2048, 30, 0),
		(drawing, 477, 7, 2048, 30, 0),
		(drawing, 478, 7, 2048, 30, 0),
		(drawing, 479, 7, 2048, 30, 0),
		(drawing, 480, 7, 2048, 30, 0),
		(drawing, 481, 7, 2048, 30, 0),
		(drawing, 482, 7, 2048, 30, 0),
		(drawing, 483, 7, 2048, 30, 0),
		(drawing, 484, 7, 2048, 30, 0),
		(drawing, 485, 7, 2048, 30, 0),
		(drawing, 486, 7, 2048, 30, 0),
		(drawing, 487, 7, 2048, 30, 0),
		(drawing, 488, 7, 2048, 30, 0),
		(drawing, 489, 7, 2048, 30, 0),
		(drawing, 490, 7, 2048, 30, 0),
		(drawing, 491, 7, 2048, 30, 0),
		(drawing, 492, 7, 2048, 30, 0),
		(drawing, 493, 7, 2048, 30, 0),
		(drawing, 494, 7, 2048, 30, 0),
		(drawing, 495, 7, 2048, 30, 0),
		(drawing, 496, 7, 2048, 30, 0),
		(drawing, 497, 7, 2048, 30, 0),
		(drawing, 498, 7, 2048, 30, 0),
		(drawing, 499, 7, 2048, 30, 0),
		(drawing, 500, 7, 2048, 30, 0),
		(drawing, 501, 7, 2048, 30, 0),
		(drawing, 502, 7, 2048, 30, 0),
		(drawing, 503, 7, 2048, 30, 0),
		(drawing, 504, 7, 2048, 30, 0),
		(drawing, 505, 7, 2048, 30, 0),
		(drawing, 506, 7, 2048, 30, 0),
		(drawing, 507, 7, 2048, 30, 0),
		(drawing, 508, 7, 2048, 30, 0),
		(drawing, 509, 7, 2048, 30, 0),
		(drawing, 510, 7, 2048, 30, 0),
		(drawing, 511, 7, 2048, 30, 0),
		(drawing, 512, 8, 2048, 30, 0),
		(drawing, 513, 8, 2048, 30, 0),
		(drawing, 514, 8, 2048, 30, 0),
		(drawing, 515, 8, 2048, 30, 0),
		(drawing, 516, 8, 2048, 30, 0),
		(drawing, 517, 8, 2048, 30, 0),
		(drawing, 518, 8, 2048, 30, 0),
		(drawing, 519, 8, 2048, 30, 0),
		(drawing, 520, 8, 2048, 30, 0),
		(drawing, 521, 8, 2048, 30, 0),
		(drawing, 522, 8, 2048, 30, 0),
		(drawing, 523, 8, 2048, 30, 0),
		(drawing, 524, 8, 2048, 30, 0),
		(drawing, 525, 8, 2048, 30, 0),
		(drawing, 526, 8, 2048, 30, 0),
		(drawing, 527, 8, 2048, 30, 0),
		(drawing, 528, 8, 2048, 30, 0),
		(drawing, 529, 8, 2048, 30, 0),
		(drawing, 530, 8, 2048, 30, 0),
		(drawing, 531, 8, 2048, 30, 0),
		(drawing, 532, 8, 2048, 30, 0),
		(drawing, 533, 8, 2048, 30, 0),
		(drawing, 534, 8, 2048, 30, 0),
		(drawing, 535, 8, 2048, 30, 0),
		(drawing, 536, 8, 2048, 30, 0),
		(drawing, 537, 8, 2048, 30, 0),
		(drawing, 538, 8, 2048, 30, 0),
		(drawing, 539, 8, 2048, 30, 0),
		(drawing, 540, 8, 2048, 30, 0),
		(drawing, 541, 8, 2048, 30, 0),
		(drawing, 542, 8, 2048, 30, 0),
		(drawing, 543, 8, 2048, 30, 0),
		(drawing, 544, 8, 2048, 30, 0),
		(drawing, 545, 8, 2048, 30, 0),
		(drawing, 546, 8, 2048, 30, 0),
		(drawing, 547, 8, 2048, 30, 0),
		(drawing, 548, 8, 2048, 30, 0),
		(drawing, 549, 8, 2048, 30, 0),
		(drawing, 550, 8, 2048, 30, 0),
		(drawing, 551, 8, 2048, 30, 0),
		(drawing, 552, 8, 2048, 30, 0),
		(drawing, 553, 8, 2048, 30, 0),
		(drawing, 554, 8, 2048, 30, 0),
		(drawing, 555, 8, 2048, 30, 0),
		(drawing, 556, 8, 2048, 30, 0),
		(drawing, 557, 8, 2048, 30, 0),
		(drawing, 558, 8, 2048, 30, 0),
		(drawing, 559, 8, 2048, 30, 0),
		(drawing, 560, 8, 2048, 30, 0),
		(drawing, 561, 8, 2048, 30, 0),
		(drawing, 562, 8, 2048, 30, 0),
		(drawing, 563, 8, 2048, 30, 0),
		(drawing, 564, 8, 2048, 30, 0),
		(drawing, 565, 8, 2048, 30, 0),
		(drawing, 566, 8, 2048, 30, 0),
		(drawing, 567, 8, 2048, 30, 0),
		(drawing, 568, 8, 2048, 30, 0),
		(drawing, 569, 8, 2048, 30, 0),
		(drawing, 570, 8, 2048, 30, 0),
		(drawing, 571, 8, 2048, 30, 0),
		(drawing, 572, 8, 2048, 30, 0),
		(drawing, 573, 8, 2048, 30, 0),
		(drawing, 574, 8, 2048, 30, 0),
		(drawing, 575, 8, 2048, 30, 0),
		(drawing, 576, 8, 2048, 30, 0),
		(drawing, 577, 8, 2048, 30, 0),
		(drawing, 578, 8, 2048, 30, 0),
		(drawing, 579, 8, 2048, 30, 0),
		(drawing, 580, 8, 2048, 30, 0),
		(drawing, 581, 9, 2048, 30, 0),
		(drawing, 582, 9, 2048, 30, 0),
		(drawing, 583, 9, 2048, 30, 0),
		(drawing, 584, 9, 2048, 30, 0),
		(drawing, 585, 9, 2048, 30, 0),
		(drawing, 586, 9, 2048, 30, 0),
		(drawing, 587, 9, 2048, 30, 0),
		(drawing, 588, 9, 2048, 30, 0),
		(drawing, 589, 9, 2048, 30, 0),
		(drawing, 590, 9, 2048, 30, 0),
		(drawing, 591, 9, 2048, 30, 0),
		(drawing, 592, 9, 2048, 30, 0),
		(drawing, 593, 9, 2048, 30, 0),
		(drawing, 594, 9, 2048, 30, 0),
		(drawing, 595, 9, 2048, 30, 0),
		(drawing, 596, 9, 2048, 30, 0),
		(drawing, 597, 9, 2048, 30, 0),
		(drawing, 598, 9, 2048, 30, 0),
		(drawing, 599, 9, 2048, 30, 0),
		(drawing, 600, 9, 2048, 30, 0),
		(drawing, 601, 9, 2048, 30, 0),
		(drawing, 602, 9, 2048, 30, 0),
		(drawing, 603, 9, 2048, 30, 0),
		(drawing, 604, 9, 2048, 30, 0),
		(drawing, 605, 9, 2048, 30, 0),
		(drawing, 606, 9, 2048, 30, 0),
		(drawing, 607, 9, 2048, 30, 0),
		(drawing, 608, 9, 2048, 30, 0),
		(drawing, 609, 9, 2048, 30, 0),
		(drawing, 610, 9, 2048, 30, 0),
		(drawing, 611, 9, 2048, 30, 0),
		(drawing, 612, 9, 2048, 30, 0),
		(drawing, 613, 9, 2048, 30, 0),
		(drawing, 614, 9, 2048, 30, 0),
		(drawing, 615, 9, 2048, 30, 0),
		(drawing, 616, 9, 2048, 30, 0),
		(drawing, 617, 9, 2048, 30, 0),
		(drawing, 618, 9, 2048, 30, 0),
		(drawing, 619, 9, 2048, 30, 0),
		(drawing, 620, 9, 2048, 30, 0),
		(drawing, 621, 9, 2048, 30, 0),
		(drawing, 622, 9, 2048, 30, 0),
		(drawing, 623, 9, 2048, 30, 0),
		(drawing, 624, 9, 2048, 30, 0),
		(drawing, 625, 9, 2048, 30, 0),
		(drawing, 626, 9, 2048, 30, 0),
		(drawing, 627, 9, 2048, 30, 0),
		(drawing, 628, 9, 2048, 30, 0),
		(drawing, 629, 9, 2048, 30, 0),
		(drawing, 630, 9, 2048, 30, 0),
		(drawing, 631, 9, 2048, 30, 0),
		(drawing, 632, 9, 2048, 30, 0),
		(drawing, 633, 9, 2048, 30, 0),
		(drawing, 634, 9, 2048, 30, 0),
		(drawing, 635, 9, 2048, 30, 0),
		(drawing, 636, 9, 2048, 30, 0),
		(drawing, 637, 9, 2048, 30, 0),
		(drawing, 638, 9, 2048, 30, 0),
		(drawing, 639, 9, 2048, 30, 0),
		(drawing, 640, 9, 2048, 30, 0),
		(drawing, 641, 9, 2048, 30, 0),
		(drawing, 642, 9, 2048, 30, 0),
		(drawing, 643, 9, 2048, 30, 0),
		(drawing, 644, 9, 2048, 30, 0),
		(drawing, 645, 9, 2048, 30, 0),
		(drawing, 646, 9, 2048, 30, 0),
		(drawing, 647, 9, 2048, 30, 0),
		(drawing, 648, 9, 2048, 30, 0),
		(drawing, 649, 10, 2048, 30, 0),
		(drawing, 650, 10, 2048, 30, 0),
		(drawing, 651, 10, 2048, 30, 0),
		(drawing, 652, 10, 2048, 30, 0),
		(drawing, 653, 10, 2048, 30, 0),
		(drawing, 654, 10, 2048, 30, 0),
		(drawing, 655, 10, 2048, 30, 0),
		(drawing, 656, 10, 2048, 30, 0),
		(drawing, 657, 10, 2048, 30, 0),
		(drawing, 658, 10, 2048, 30, 0),
		(drawing, 659, 10, 2048, 30, 0),
		(drawing, 660, 10, 2048, 30, 0),
		(drawing, 661, 10, 2048, 30, 0),
		(drawing, 662, 10, 2048, 30, 0),
		(drawing, 663, 10, 2048, 30, 0),
		(drawing, 664, 10, 2048, 30, 0),
		(drawing, 665, 10, 2048, 30, 0),
		(drawing, 666, 10, 2048, 30, 0),
		(drawing, 667, 10, 2048, 30, 0),
		(drawing, 668, 10, 2048, 30, 0),
		(drawing, 669, 10, 2048, 30, 0),
		(drawing, 670, 10, 2048, 30, 0),
		(drawing, 671, 10, 2048, 30, 0),
		(drawing, 672, 10, 2048, 30, 0),
		(drawing, 673, 10, 2048, 30, 0),
		(drawing, 674, 10, 2048, 30, 0),
		(drawing, 675, 10, 2048, 30, 0),
		(drawing, 676, 10, 2048, 30, 0),
		(drawing, 677, 10, 2048, 30, 0),
		(drawing, 678, 10, 2048, 30, 0),
		(drawing, 679, 10, 2048, 30, 0),
		(drawing, 680, 10, 2048, 30, 0),
		(drawing, 681, 10, 2048, 30, 0),
		(drawing, 682, 10, 2048, 30, 0),
		(drawing, 683, 10, 2048, 30, 0),
		(drawing, 684, 10, 2048, 30, 0),
		(drawing, 685, 10, 2048, 30, 0),
		(drawing, 686, 10, 2048, 30, 0),
		(drawing, 687, 10, 2048, 30, 0),
		(drawing, 688, 10, 2048, 30, 0),
		(drawing, 689, 10, 2048, 30, 0),
		(drawing, 690, 10, 2048, 30, 0),
		(drawing, 691, 10, 2048, 30, 0),
		(drawing, 692, 10, 2048, 30, 0),
		(drawing, 693, 10, 2048, 30, 0),
		(drawing, 694, 10, 2048, 30, 0),
		(drawing, 695, 10, 2048, 30, 0),
		(drawing, 696, 10, 2048, 30, 0),
		(drawing, 697, 10, 2048, 30, 0),
		(drawing, 698, 10, 2048, 30, 0),
		(drawing, 699, 10, 2048, 30, 0),
		(drawing, 700, 10, 2048, 30, 0),
		(drawing, 701, 10, 2048, 30, 0),
		(drawing, 702, 10, 2048, 30, 0),
		(drawing, 703, 10, 2048, 30, 0),
		(drawing, 704, 10, 2048, 30, 0),
		(drawing, 705, 10, 2048, 30, 0),
		(drawing, 706, 10, 2048, 30, 0),
		(drawing, 707, 10, 2048, 30, 0),
		(drawing, 708, 10, 2048, 30, 0),
		(drawing, 709, 10, 2048, 30, 0),
		(drawing, 710, 10, 2048, 30, 0),
		(drawing, 711, 10, 2048, 30, 0),
		(drawing, 712, 10, 2048, 30, 0),
		(drawing, 713, 10, 2048, 30, 0),
		(drawing, 714, 10, 2048, 30, 0),
		(drawing, 715, 10, 2048, 30, 0),
		(drawing, 716, 10, 2048, 30, 0),
		(drawing, 717, 11, 2048, 30, 0),
		(drawing, 718, 11, 2048, 30, 0),
		(drawing, 719, 11, 2048, 30, 0),
		(drawing, 720, 11, 2048, 30, 0),
		(drawing, 721, 11, 2048, 30, 0),
		(drawing, 722, 11, 2048, 30, 0),
		(drawing, 723, 11, 2048, 30, 0),
		(drawing, 724, 11, 2048, 30, 0),
		(drawing, 725, 11, 2048, 30, 0),
		(drawing, 726, 11, 2048, 30, 0),
		(drawing, 727, 11, 2048, 30, 0),
		(drawing, 728, 11, 2048, 30, 0),
		(drawing, 729, 11, 2048, 30, 0),
		(drawing, 730, 11, 2048, 30, 0),
		(drawing, 731, 11, 2048, 30, 0),
		(drawing, 732, 11, 2048, 30, 0),
		(drawing, 733, 11, 2048, 30, 0),
		(drawing, 734, 11, 2048, 30, 0),
		(drawing, 735, 11, 2048, 30, 0),
		(drawing, 736, 11, 2048, 30, 0),
		(drawing, 737, 11, 2048, 30, 0),
		(drawing, 738, 11, 2048, 30, 0),
		(drawing, 739, 11, 2048, 30, 0),
		(drawing, 740, 11, 2048, 30, 0),
		(drawing, 741, 11, 2048, 30, 0),
		(drawing, 742, 11, 2048, 30, 0),
		(drawing, 743, 11, 2048, 30, 0),
		(drawing, 744, 11, 2048, 30, 0),
		(drawing, 745, 11, 2048, 30, 0),
		(drawing, 746, 11, 2048, 30, 0),
		(drawing, 747, 11, 2048, 30, 0),
		(drawing, 748, 11, 2048, 30, 0),
		(drawing, 749, 11, 2048, 30, 0),
		(drawing, 750, 11, 2048, 30, 0),
		(drawing, 751, 11, 2048, 30, 0),
		(drawing, 752, 11, 2048, 30, 0),
		(drawing, 753, 11, 2048, 30, 0),
		(drawing, 754, 11, 2048, 30, 0),
		(drawing, 755, 11, 2048, 30, 0),
		(drawing, 756, 11, 2048, 30, 0),
		(drawing, 757, 11, 2048, 30, 0),
		(drawing, 758, 11, 2048, 30, 0),
		(drawing, 759, 11, 2048, 30, 0),
		(drawing, 760, 11, 2048, 30, 0),
		(drawing, 761, 11, 2048, 30, 0),
		(drawing, 762, 11, 2048, 30, 0),
		(drawing, 763, 11, 2048, 30, 0),
		(drawing, 764, 11, 2048, 30, 0),
		(drawing, 765, 11, 2048, 30, 0),
		(drawing, 766, 11, 2048, 30, 0),
		(drawing, 767, 11, 2048, 30, 0),
		(drawing, 768, 11, 2048, 30, 0),
		(drawing, 769, 11, 2048, 30, 0),
		(drawing, 770, 11, 2048, 30, 0),
		(drawing, 771, 11, 2048, 30, 0),
		(drawing, 772, 11, 2048, 30, 0),
		(drawing, 773, 11, 2048, 30, 0),
		(drawing, 774, 11, 2048, 30, 0),
		(drawing, 775, 11, 2048, 30, 0),
		(drawing, 776, 11, 2048, 30, 0),
		(drawing, 777, 11, 2048, 30, 0),
		(drawing, 778, 11, 2048, 30, 0),
		(drawing, 779, 11, 2048, 30, 0),
		(drawing, 780, 11, 2048, 30, 0),
		(drawing, 781, 11, 2048, 30, 0),
		(drawing, 782, 11, 2048, 30, 0),
		(drawing, 783, 11, 2048, 30, 0),
		(drawing, 784, 11, 2048, 30, 0),
		(drawing, 785, 11, 2048, 30, 0),
		(drawing, 786, 12, 2048, 30, 0),
		(drawing, 787, 12, 2048, 30, 0),
		(drawing, 788, 12, 2048, 30, 0),
		(drawing, 789, 12, 2048, 30, 0),
		(drawing, 790, 12, 2048, 30, 0),
		(drawing, 791, 12, 2048, 30, 0),
		(drawing, 792, 12, 2048, 30, 0),
		(drawing, 793, 12, 2048, 30, 0),
		(drawing, 794, 12, 2048, 30, 0),
		(drawing, 795, 12, 2048, 30, 0),
		(drawing, 796, 12, 2048, 30, 0),
		(drawing, 797, 12, 2048, 30, 0),
		(drawing, 798, 12, 2048, 30, 0),
		(drawing, 799, 12, 2048, 30, 0),
		(drawing, 800, 12, 2048, 30, 0),
		(drawing, 801, 12, 2048, 30, 0),
		(drawing, 802, 12, 2048, 30, 0),
		(drawing, 803, 12, 2048, 30, 0),
		(drawing, 804, 12, 2048, 30, 0),
		(drawing, 805, 12, 2048, 30, 0),
		(drawing, 806, 12, 2048, 30, 0),
		(drawing, 807, 12, 2048, 30, 0),
		(drawing, 808, 12, 2048, 30, 0),
		(drawing, 809, 12, 2048, 30, 0),
		(drawing, 810, 12, 2048, 30, 0),
		(drawing, 811, 12, 2048, 30, 0),
		(drawing, 812, 12, 2048, 30, 0),
		(drawing, 813, 12, 2048, 30, 0),
		(drawing, 814, 12, 2048, 30, 0),
		(drawing, 815, 12, 2048, 30, 0),
		(drawing, 816, 12, 2048, 30, 0),
		(drawing, 817, 12, 2048, 30, 0),
		(drawing, 818, 12, 2048, 30, 0),
		(drawing, 819, 12, 2048, 30, 0),
		(drawing, 820, 12, 2048, 30, 0),
		(drawing, 821, 12, 2048, 30, 0),
		(drawing, 822, 12, 2048, 30, 0),
		(drawing, 823, 12, 2048, 30, 0),
		(drawing, 824, 12, 2048, 30, 0),
		(drawing, 825, 12, 2048, 30, 0),
		(drawing, 826, 12, 2048, 30, 0),
		(drawing, 827, 12, 2048, 30, 0),
		(drawing, 828, 12, 2048, 30, 0),
		(drawing, 829, 12, 2048, 30, 0),
		(drawing, 830, 12, 2048, 30, 0),
		(drawing, 831, 12, 2048, 30, 0),
		(drawing, 832, 12, 2048, 30, 0),
		(drawing, 833, 12, 2048, 30, 0),
		(drawing, 834, 12, 2048, 30, 0),
		(drawing, 835, 12, 2048, 30, 0),
		(drawing, 836, 12, 2048, 30, 0),
		(drawing, 837, 12, 2048, 30, 0),
		(drawing, 838, 12, 2048, 30, 0),
		(drawing, 839, 12, 2048, 30, 0),
		(drawing, 840, 12, 2048, 30, 0),
		(drawing, 841, 12, 2048, 30, 0),
		(drawing, 842, 12, 2048, 30, 0),
		(drawing, 843, 12, 2048, 30, 0),
		(drawing, 844, 12, 2048, 30, 0),
		(drawing, 845, 12, 2048, 30, 0),
		(drawing, 846, 12, 2048, 30, 0),
		(drawing, 847, 12, 2048, 30, 0),
		(drawing, 848, 12, 2048, 30, 0),
		(drawing, 849, 12, 2048, 30, 0),
		(drawing, 850, 12, 2048, 30, 0),
		(drawing, 851, 12, 2048, 30, 0),
		(drawing, 852, 12, 2048, 30, 0),
		(drawing, 853, 12, 2048, 30, 0),
		(drawing, 854, 13, 2048, 30, 0),
		(drawing, 855, 13, 2048, 30, 0),
		(drawing, 856, 13, 2048, 30, 0),
		(drawing, 857, 13, 2048, 30, 0),
		(drawing, 858, 13, 2048, 30, 0),
		(drawing, 859, 13, 2048, 30, 0),
		(drawing, 860, 13, 2048, 30, 0),
		(drawing, 861, 13, 2048, 30, 0),
		(drawing, 862, 13, 2048, 30, 0),
		(drawing, 863, 13, 2048, 30, 0),
		(drawing, 864, 13, 2048, 30, 0),
		(drawing, 865, 13, 2048, 30, 0),
		(drawing, 866, 13, 2048, 30, 0),
		(drawing, 867, 13, 2048, 30, 0),
		(drawing, 868, 13, 2048, 30, 0),
		(drawing, 869, 13, 2048, 30, 0),
		(drawing, 870, 13, 2048, 30, 0),
		(drawing, 871, 13, 2048, 30, 0),
		(drawing, 872, 13, 2048, 30, 0),
		(drawing, 873, 13, 2048, 30, 0),
		(drawing, 874, 13, 2048, 30, 0),
		(drawing, 875, 13, 2048, 30, 0),
		(drawing, 876, 13, 2048, 30, 0),
		(drawing, 877, 13, 2048, 30, 0),
		(drawing, 878, 13, 2048, 30, 0),
		(drawing, 879, 13, 2048, 30, 0),
		(drawing, 880, 13, 2048, 30, 0),
		(drawing, 881, 13, 2048, 30, 0),
		(drawing, 882, 13, 2048, 30, 0),
		(drawing, 883, 13, 2048, 30, 0),
		(drawing, 884, 13, 2048, 30, 0),
		(drawing, 885, 13, 2048, 30, 0),
		(drawing, 886, 13, 2048, 30, 0),
		(drawing, 887, 13, 2048, 30, 0),
		(drawing, 888, 13, 2048, 30, 0),
		(drawing, 889, 13, 2048, 30, 0),
		(drawing, 890, 13, 2048, 30, 0),
		(drawing, 891, 13, 2048, 30, 0),
		(drawing, 892, 13, 2048, 30, 0),
		(drawing, 893, 13, 2048, 30, 0),
		(drawing, 894, 13, 2048, 30, 0),
		(drawing, 895, 13, 2048, 30, 0),
		(drawing, 896, 13, 2048, 30, 0),
		(drawing, 897, 13, 2048, 30, 0),
		(drawing, 898, 13, 2048, 30, 0),
		(drawing, 899, 13, 2048, 30, 0),
		(drawing, 900, 13, 2048, 30, 0),
		(drawing, 901, 13, 2048, 30, 0),
		(drawing, 902, 13, 2048, 30, 0),
		(drawing, 903, 13, 2048, 30, 0),
		(drawing, 904, 13, 2048, 30, 0),
		(drawing, 905, 13, 2048, 30, 0),
		(drawing, 906, 13, 2048, 30, 0),
		(drawing, 907, 13, 2048, 30, 0),
		(drawing, 908, 13, 2048, 30, 0),
		(drawing, 909, 13, 2048, 30, 0),
		(drawing, 910, 13, 2048, 30, 0),
		(drawing, 911, 13, 2048, 30, 0),
		(drawing, 912, 13, 2048, 30, 0),
		(drawing, 913, 13, 2048, 30, 0),
		(drawing, 914, 13, 2048, 30, 0),
		(drawing, 915, 13, 2048, 30, 0),
		(drawing, 916, 13, 2048, 30, 0),
		(drawing, 917, 13, 2048, 30, 0),
		(drawing, 918, 13, 2048, 30, 0),
		(drawing, 919, 13, 2048, 30, 0),
		(drawing, 920, 13, 2048, 30, 0),
		(drawing, 921, 13, 2048, 30, 0),
		(drawing, 922, 14, 2048, 30, 0),
		(drawing, 923, 14, 2048, 30, 0),
		(drawing, 924, 14, 2048, 30, 0),
		(drawing, 925, 14, 2048, 30, 0),
		(drawing, 926, 14, 2048, 30, 0),
		(drawing, 927, 14, 2048, 30, 0),
		(drawing, 928, 14, 2048, 30, 0),
		(drawing, 929, 14, 2048, 30, 0),
		(drawing, 930, 14, 2048, 30, 0),
		(drawing, 931, 14, 2048, 30, 0),
		(drawing, 932, 14, 2048, 30, 0),
		(drawing, 933, 14, 2048, 30, 0),
		(drawing, 934, 14, 2048, 30, 0),
		(drawing, 935, 14, 2048, 30, 0),
		(drawing, 936, 14, 2048, 30, 0),
		(drawing, 937, 14, 2048, 30, 0),
		(drawing, 938, 14, 2048, 30, 0),
		(drawing, 939, 14, 2048, 30, 0),
		(drawing, 940, 14, 2048, 30, 0),
		(drawing, 941, 14, 2048, 30, 0),
		(drawing, 942, 14, 2048, 30, 0),
		(drawing, 943, 14, 2048, 30, 0),
		(drawing, 944, 14, 2048, 30, 0),
		(drawing, 945, 14, 2048, 30, 0),
		(drawing, 946, 14, 2048, 30, 0),
		(drawing, 947, 14, 2048, 30, 0),
		(drawing, 948, 14, 2048, 30, 0),
		(drawing, 949, 14, 2048, 30, 0),
		(drawing, 950, 14, 2048, 30, 0),
		(drawing, 951, 14, 2048, 30, 0),
		(drawing, 952, 14, 2048, 30, 0),
		(drawing, 953, 14, 2048, 30, 0),
		(drawing, 954, 14, 2048, 30, 0),
		(drawing, 955, 14, 2048, 30, 0),
		(drawing, 956, 14, 2048, 30, 0),
		(drawing, 957, 14, 2048, 30, 0),
		(drawing, 958, 14, 2048, 30, 0),
		(drawing, 959, 14, 2048, 30, 0),
		(drawing, 960, 14, 2048, 30, 0),
		(drawing, 961, 14, 2048, 30, 0),
		(drawing, 962, 14, 2048, 30, 0),
		(drawing, 963, 14, 2048, 30, 0),
		(drawing, 964, 14, 2048, 30, 0),
		(drawing, 965, 14, 2048, 30, 0),
		(drawing, 966, 14, 2048, 30, 0),
		(drawing, 967, 14, 2048, 30, 0),
		(drawing, 968, 14, 2048, 30, 0),
		(drawing, 969, 14, 2048, 30, 0),
		(drawing, 970, 14, 2048, 30, 0),
		(drawing, 971, 14, 2048, 30, 0),
		(drawing, 972, 14, 2048, 30, 0),
		(drawing, 973, 14, 2048, 30, 0),
		(drawing, 974, 14, 2048, 30, 0),
		(drawing, 975, 14, 2048, 30, 0),
		(drawing, 976, 14, 2048, 30, 0),
		(drawing, 977, 14, 2048, 30, 0),
		(drawing, 978, 14, 2048, 30, 0),
		(drawing, 979, 14, 2048, 30, 0),
		(drawing, 980, 14, 2048, 30, 0),
		(drawing, 981, 14, 2048, 30, 0),
		(drawing, 982, 14, 2048, 30, 0),
		(drawing, 983, 14, 2048, 30, 0),
		(drawing, 984, 14, 2048, 30, 0),
		(drawing, 985, 14, 2048, 30, 0),
		(drawing, 986, 14, 2048, 30, 0),
		(drawing, 987, 14, 2048, 30, 0),
		(drawing, 988, 14, 2048, 30, 0),
		(drawing, 989, 14, 2048, 30, 0),
		(drawing, 990, 15, 2048, 30, 0),
		(drawing, 991, 15, 2048, 30, 0),
		(drawing, 992, 15, 2048, 30, 0),
		(drawing, 993, 15, 2048, 30, 0),
		(drawing, 994, 15, 2048, 30, 0),
		(drawing, 995, 15, 2048, 30, 0),
		(drawing, 996, 15, 2048, 30, 0),
		(drawing, 997, 15, 2048, 30, 0),
		(drawing, 998, 15, 2048, 30, 0),
		(drawing, 999, 15, 2048, 30, 0),
		(drawing, 1000, 15, 2048, 30, 0),
		(drawing, 1001, 15, 2048, 30, 0),
		(drawing, 1002, 15, 2048, 30, 0),
		(drawing, 1003, 15, 2048, 30, 0),
		(drawing, 1004, 15, 2048, 30, 0),
		(drawing, 1005, 15, 2048, 30, 0),
		(drawing, 1006, 15, 2048, 30, 0),
		(drawing, 1007, 15, 2048, 30, 0),
		(drawing, 1008, 15, 2048, 30, 0),
		(drawing, 1009, 15, 2048, 30, 0),
		(drawing, 1010, 15, 2048, 30, 0),
		(drawing, 1011, 15, 2048, 30, 0),
		(drawing, 1012, 15, 2048, 30, 0),
		(drawing, 1013, 15, 2048, 30, 0),
		(drawing, 1014, 15, 2048, 30, 0),
		(drawing, 1015, 15, 2048, 30, 0),
		(drawing, 1016, 15, 2048, 30, 0),
		(drawing, 1017, 15, 2048, 30, 0),
		(drawing, 1018, 15, 2048, 30, 0),
		(drawing, 1019, 15, 2048, 30, 0),
		(drawing, 1020, 15, 2048, 30, 0),
		(drawing, 1021, 15, 2048, 30, 0),
		(drawing, 1022, 15, 2048, 30, 0),
		(drawing, 1023, 15, 2048, 30, 0),
		(drawing, 1024, 15, 2048, 30, 0),
		(drawing, 1025, 15, 2048, 30, 0),
		(drawing, 1026, 15, 2048, 30, 0),
		(drawing, 1027, 15, 2048, 30, 0),
		(drawing, 1028, 15, 2048, 30, 0),
		(drawing, 1029, 15, 2048, 30, 0),
		(drawing, 1030, 15, 2048, 30, 0),
		(drawing, 1031, 15, 2048, 30, 0),
		(drawing, 1032, 15, 2048, 30, 0),
		(drawing, 1033, 15, 2048, 30, 0),
		(drawing, 1034, 15, 2048, 30, 0),
		(drawing, 1035, 15, 2048, 30, 0),
		(drawing, 1036, 15, 2048, 30, 0),
		(drawing, 1037, 15, 2048, 30, 0),
		(drawing, 1038, 15, 2048, 30, 0),
		(drawing, 1039, 15, 2048, 30, 0),
		(drawing, 1040, 15, 2048, 30, 0),
		(drawing, 1041, 15, 2048, 30, 0),
		(drawing, 1042, 15, 2048, 30, 0),
		(drawing, 1043, 15, 2048, 30, 0),
		(drawing, 1044, 15, 2048, 30, 0),
		(drawing, 1045, 15, 2048, 30, 0),
		(drawing, 1046, 15, 2048, 30, 0),
		(drawing, 1047, 15, 2048, 30, 0),
		(drawing, 1048, 15, 2048, 30, 0),
		(drawing, 1049, 15, 2048, 30, 0),
		(drawing, 1050, 15, 2048, 30, 0),
		(drawing, 1051, 15, 2048, 30, 0),
		(drawing, 1052, 15, 2048, 30, 0),
		(drawing, 1053, 15, 2048, 30, 0),
		(drawing, 1054, 15, 2048, 30, 0),
		(drawing, 1055, 15, 2048, 30, 0),
		(drawing, 1056, 15, 2048, 30, 0),
		(drawing, 1057, 15, 2048, 30, 0),
		(drawing, 1058, 15, 2048, 30, 0),
		(drawing, 1059, 16, 2048, 30, 0),
		(drawing, 1060, 16, 2048, 30, 0),
		(drawing, 1061, 16, 2048, 30, 0),
		(drawing, 1062, 16, 2048, 30, 0),
		(drawing, 1063, 16, 2048, 30, 0),
		(drawing, 1064, 16, 2048, 30, 0),
		(drawing, 1065, 16, 2048, 30, 0),
		(drawing, 1066, 16, 2048, 30, 0),
		(drawing, 1067, 16, 2048, 30, 0),
		(drawing, 1068, 16, 2048, 30, 0),
		(drawing, 1069, 16, 2048, 30, 0),
		(drawing, 1070, 16, 2048, 30, 0),
		(drawing, 1071, 16, 2048, 30, 0),
		(drawing, 1072, 16, 2048, 30, 0),
		(drawing, 1073, 16, 2048, 30, 0),
		(drawing, 1074, 16, 2048, 30, 0),
		(drawing, 1075, 16, 2048, 30, 0),
		(drawing, 1076, 16, 2048, 30, 0),
		(drawing, 1077, 16, 2048, 30, 0),
		(drawing, 1078, 16, 2048, 30, 0),
		(drawing, 1079, 16, 2048, 30, 0),
		(drawing, 1080, 16, 2048, 30, 0),
		(drawing, 1081, 16, 2048, 30, 0),
		(drawing, 1082, 16, 2048, 30, 0),
		(drawing, 1083, 16, 2048, 30, 0),
		(drawing, 1084, 16, 2048, 30, 0),
		(drawing, 1085, 16, 2048, 30, 0),
		(drawing, 1086, 16, 2048, 30, 0),
		(drawing, 1087, 16, 2048, 30, 0),
		(drawing, 1088, 16, 2048, 30, 0),
		(drawing, 1089, 16, 2048, 30, 0),
		(drawing, 1090, 16, 2048, 30, 0),
		(drawing, 1091, 16, 2048, 30, 0),
		(drawing, 1092, 16, 2048, 30, 0),
		(drawing, 1093, 16, 2048, 30, 0),
		(drawing, 1094, 16, 2048, 30, 0),
		(drawing, 1095, 16, 2048, 30, 0),
		(drawing, 1096, 16, 2048, 30, 0),
		(drawing, 1097, 16, 2048, 30, 0),
		(drawing, 1098, 16, 2048, 30, 0),
		(drawing, 1099, 16, 2048, 30, 0),
		(drawing, 1100, 16, 2048, 30, 0),
		(drawing, 1101, 16, 2048, 30, 0),
		(drawing, 1102, 16, 2048, 30, 0),
		(drawing, 1103, 16, 2048, 30, 0),
		(drawing, 1104, 16, 2048, 30, 0),
		(drawing, 1105, 16, 2048, 30, 0),
		(drawing, 1106, 16, 2048, 30, 0),
		(drawing, 1107, 16, 2048, 30, 0),
		(drawing, 1108, 16, 2048, 30, 0),
		(drawing, 1109, 16, 2048, 30, 0),
		(drawing, 1110, 16, 2048, 30, 0),
		(drawing, 1111, 16, 2048, 30, 0),
		(drawing, 1112, 16, 2048, 30, 0),
		(drawing, 1113, 16, 2048, 30, 0),
		(drawing, 1114, 16, 2048, 30, 0),
		(drawing, 1115, 16, 2048, 30, 0),
		(drawing, 1116, 16, 2048, 30, 0),
		(drawing, 1117, 16, 2048, 30, 0),
		(drawing, 1118, 16, 2048, 30, 0),
		(drawing, 1119, 16, 2048, 30, 0),
		(drawing, 1120, 16, 2048, 30, 0),
		(drawing, 1121, 16, 2048, 30, 0),
		(drawing, 1122, 16, 2048, 30, 0),
		(drawing, 1123, 16, 2048, 30, 0),
		(drawing, 1124, 16, 2048, 30, 0),
		(drawing, 1125, 16, 2048, 30, 0),
		(drawing, 1126, 16, 2048, 30, 0),
		(drawing, 1127, 17, 2048, 30, 0),
		(drawing, 1128, 17, 2048, 30, 0),
		(drawing, 1129, 17, 2048, 30, 0),
		(drawing, 1130, 17, 2048, 30, 0),
		(drawing, 1131, 17, 2048, 30, 0),
		(drawing, 1132, 17, 2048, 30, 0),
		(drawing, 1133, 17, 2048, 30, 0),
		(drawing, 1134, 17, 2048, 30, 0),
		(drawing, 1135, 17, 2048, 30, 0),
		(drawing, 1136, 17, 2048, 30, 0),
		(drawing, 1137, 17, 2048, 30, 0),
		(drawing, 1138, 17, 2048, 30, 0),
		(drawing, 1139, 17, 2048, 30, 0),
		(drawing, 1140, 17, 2048, 30, 0),
		(drawing, 1141, 17, 2048, 30, 0),
		(drawing, 1142, 17, 2048, 30, 0),
		(drawing, 1143, 17, 2048, 30, 0),
		(drawing, 1144, 17, 2048, 30, 0),
		(drawing, 1145, 17, 2048, 30, 0),
		(drawing, 1146, 17, 2048, 30, 0),
		(drawing, 1147, 17, 2048, 30, 0),
		(drawing, 1148, 17, 2048, 30, 0),
		(drawing, 1149, 17, 2048, 30, 0),
		(drawing, 1150, 17, 2048, 30, 0),
		(drawing, 1151, 17, 2048, 30, 0),
		(drawing, 1152, 17, 2048, 30, 0),
		(drawing, 1153, 17, 2048, 30, 0),
		(drawing, 1154, 17, 2048, 30, 0),
		(drawing, 1155, 17, 2048, 30, 0),
		(drawing, 1156, 17, 2048, 30, 0),
		(drawing, 1157, 17, 2048, 30, 0),
		(drawing, 1158, 17, 2048, 30, 0),
		(drawing, 1159, 17, 2048, 30, 0),
		(drawing, 1160, 17, 2048, 30, 0),
		(drawing, 1161, 17, 2048, 30, 0),
		(drawing, 1162, 17, 2048, 30, 0),
		(drawing, 1163, 17, 2048, 30, 0),
		(drawing, 1164, 17, 2048, 30, 0),
		(drawing, 1165, 17, 2048, 30, 0),
		(drawing, 1166, 17, 2048, 30, 0),
		(drawing, 1167, 17, 2048, 30, 0),
		(drawing, 1168, 17, 2048, 30, 0),
		(drawing, 1169, 17, 2048, 30, 0),
		(drawing, 1170, 17, 2048, 30, 0),
		(drawing, 1171, 17, 2048, 30, 0),
		(drawing, 1172, 17, 2048, 30, 0),
		(drawing, 1173, 17, 2048, 30, 0),
		(drawing, 1174, 17, 2048, 30, 0),
		(drawing, 1175, 17, 2048, 30, 0),
		(drawing, 1176, 17, 2048, 30, 0),
		(drawing, 1177, 17, 2048, 30, 0),
		(drawing, 1178, 17, 2048, 30, 0),
		(drawing, 1179, 17, 2048, 30, 0),
		(drawing, 1180, 17, 2048, 30, 0),
		(drawing, 1181, 17, 2048, 30, 0),
		(drawing, 1182, 17, 2048, 30, 0),
		(drawing, 1183, 17, 2048, 30, 0),
		(drawing, 1184, 17, 2048, 30, 0),
		(drawing, 1185, 17, 2048, 30, 0),
		(drawing, 1186, 17, 2048, 30, 0),
		(drawing, 1187, 17, 2048, 30, 0),
		(drawing, 1188, 17, 2048, 30, 0),
		(drawing, 1189, 17, 2048, 30, 0),
		(drawing, 1190, 17, 2048, 30, 0),
		(drawing, 1191, 17, 2048, 30, 0),
		(drawing, 1192, 17, 2048, 30, 0),
		(drawing, 1193, 17, 2048, 30, 0),
		(drawing, 1194, 17, 2048, 30, 0),
		(drawing, 1195, 18, 2048, 30, 0),
		(drawing, 1196, 18, 2048, 30, 0),
		(drawing, 1197, 18, 2048, 30, 0),
		(drawing, 1198, 18, 2048, 30, 0),
		(drawing, 1199, 18, 2048, 30, 0),
		(drawing, 1200, 18, 2048, 30, 0),
		(drawing, 1201, 18, 2048, 30, 0),
		(drawing, 1202, 18, 2048, 30, 0),
		(drawing, 1203, 18, 2048, 30, 0),
		(drawing, 1204, 18, 2048, 30, 0),
		(drawing, 1205, 18, 2048, 30, 0),
		(drawing, 1206, 18, 2048, 30, 0),
		(drawing, 1207, 18, 2048, 30, 0),
		(drawing, 1208, 18, 2048, 30, 0),
		(drawing, 1209, 18, 2048, 30, 0),
		(drawing, 1210, 18, 2048, 30, 0),
		(drawing, 1211, 18, 2048, 30, 0),
		(drawing, 1212, 18, 2048, 30, 0),
		(drawing, 1213, 18, 2048, 30, 0),
		(drawing, 1214, 18, 2048, 30, 0),
		(drawing, 1215, 18, 2048, 30, 0),
		(drawing, 1216, 18, 2048, 30, 0),
		(drawing, 1217, 18, 2048, 30, 0),
		(drawing, 1218, 18, 2048, 30, 0),
		(drawing, 1219, 18, 2048, 30, 0),
		(drawing, 1220, 18, 2048, 30, 0),
		(drawing, 1221, 18, 2048, 30, 0),
		(drawing, 1222, 18, 2048, 30, 0),
		(drawing, 1223, 18, 2048, 30, 0),
		(drawing, 1224, 18, 2048, 30, 0),
		(drawing, 1225, 18, 2048, 30, 0),
		(drawing, 1226, 18, 2048, 30, 0),
		(drawing, 1227, 18, 2048, 30, 0),
		(drawing, 1228, 18, 2048, 30, 0),
		(drawing, 1229, 18, 2048, 30, 0),
		(drawing, 1230, 18, 2048, 30, 0),
		(drawing, 1231, 18, 2048, 30, 0),
		(drawing, 1232, 18, 2048, 30, 0),
		(drawing, 1233, 18, 2048, 30, 0),
		(drawing, 1234, 18, 2048, 30, 0),
		(drawing, 1235, 18, 2048, 30, 0),
		(drawing, 1236, 18, 2048, 30, 0),
		(drawing, 1237, 18, 2048, 30, 0),
		(drawing, 1238, 18, 2048, 30, 0),
		(drawing, 1239, 18, 2048, 30, 0),
		(drawing, 1240, 18, 2048, 30, 0),
		(drawing, 1241, 18, 2048, 30, 0),
		(drawing, 1242, 18, 2048, 30, 0),
		(drawing, 1243, 18, 2048, 30, 0),
		(drawing, 1244, 18, 2048, 30, 0),
		(drawing, 1245, 18, 2048, 30, 0),
		(drawing, 1246, 18, 2048, 30, 0),
		(drawing, 1247, 18, 2048, 30, 0),
		(drawing, 1248, 18, 2048, 30, 0),
		(drawing, 1249, 18, 2048, 30, 0),
		(drawing, 1250, 18, 2048, 30, 0),
		(drawing, 1251, 18, 2048, 30, 0),
		(drawing, 1252, 18, 2048, 30, 0),
		(drawing, 1253, 18, 2048, 30, 0),
		(drawing, 1254, 18, 2048, 30, 0),
		(drawing, 1255, 18, 2048, 30, 0),
		(drawing, 1256, 18, 2048, 30, 0),
		(drawing, 1257, 18, 2048, 30, 0),
		(drawing, 1258, 18, 2048, 30, 0),
		(drawing, 1259, 18, 2048, 30, 0),
		(drawing, 1260, 18, 2048, 30, 0),
		(drawing, 1261, 18, 2048, 30, 0),
		(drawing, 1262, 18, 2048, 30, 0),
		(drawing, 1263, 19, 2048, 30, 0),
		(drawing, 1264, 19, 2048, 30, 0),
		(drawing, 1265, 19, 2048, 30, 0),
		(drawing, 1266, 19, 2048, 30, 0),
		(drawing, 1267, 19, 2048, 30, 0),
		(drawing, 1268, 19, 2048, 30, 0),
		(drawing, 1269, 19, 2048, 30, 0),
		(drawing, 1270, 19, 2048, 30, 0),
		(drawing, 1271, 19, 2048, 30, 0),
		(drawing, 1272, 19, 2048, 30, 0),
		(drawing, 1273, 19, 2048, 30, 0),
		(drawing, 1274, 19, 2048, 30, 0),
		(drawing, 1275, 19, 2048, 30, 0),
		(drawing, 1276, 19, 2048, 30, 0),
		(drawing, 1277, 19, 2048, 30, 0),
		(drawing, 1278, 19, 2048, 30, 0),
		(drawing, 1279, 19, 2048, 30, 0),
		(drawing, 1280, 19, 2048, 30, 0),
		(drawing, 1281, 19, 2048, 30, 0),
		(drawing, 1282, 19, 2048, 30, 0),
		(drawing, 1283, 19, 2048, 30, 0),
		(drawing, 1284, 19, 2048, 30, 0),
		(drawing, 1285, 19, 2048, 30, 0),
		(drawing, 1286, 19, 2048, 30, 0),
		(drawing, 1287, 19, 2048, 30, 0),
		(drawing, 1288, 19, 2048, 30, 0),
		(drawing, 1289, 19, 2048, 30, 0),
		(drawing, 1290, 19, 2048, 30, 0),
		(drawing, 1291, 19, 2048, 30, 0),
		(drawing, 1292, 19, 2048, 30, 0),
		(drawing, 1293, 19, 2048, 30, 0),
		(drawing, 1294, 19, 2048, 30, 0),
		(drawing, 1295, 19, 2048, 30, 0),
		(drawing, 1296, 19, 2048, 30, 0),
		(drawing, 1297, 19, 2048, 30, 0),
		(drawing, 1298, 19, 2048, 30, 0),
		(drawing, 1299, 19, 2048, 30, 0),
		(drawing, 1300, 19, 2048, 30, 0),
		(drawing, 1301, 19, 2048, 30, 0),
		(drawing, 1302, 19, 2048, 30, 0),
		(drawing, 1303, 19, 2048, 30, 0),
		(drawing, 1304, 19, 2048, 30, 0),
		(drawing, 1305, 19, 2048, 30, 0),
		(drawing, 1306, 19, 2048, 30, 0),
		(drawing, 1307, 19, 2048, 30, 0),
		(drawing, 1308, 19, 2048, 30, 0),
		(drawing, 1309, 19, 2048, 30, 0),
		(drawing, 1310, 19, 2048, 30, 0),
		(drawing, 1311, 19, 2048, 30, 0),
		(drawing, 1312, 19, 2048, 30, 0),
		(drawing, 1313, 19, 2048, 30, 0),
		(drawing, 1314, 19, 2048, 30, 0),
		(drawing, 1315, 19, 2048, 30, 0),
		(drawing, 1316, 19, 2048, 30, 0),
		(drawing, 1317, 19, 2048, 30, 0),
		(drawing, 1318, 19, 2048, 30, 0),
		(drawing, 1319, 19, 2048, 30, 0),
		(drawing, 1320, 19, 2048, 30, 0),
		(drawing, 1321, 19, 2048, 30, 0),
		(drawing, 1322, 19, 2048, 30, 0),
		(drawing, 1323, 19, 2048, 30, 0),
		(drawing, 1324, 19, 2048, 30, 0),
		(drawing, 1325, 19, 2048, 30, 0),
		(drawing, 1326, 19, 2048, 30, 0),
		(drawing, 1327, 19, 2048, 30, 0),
		(drawing, 1328, 19, 2048, 30, 0),
		(drawing, 1329, 19, 2048, 30, 0),
		(drawing, 1330, 19, 2048, 30, 0),
		(drawing, 1331, 19, 2048, 30, 0),
		(drawing, 1332, 20, 2048, 30, 0),
		(drawing, 1333, 20, 2048, 30, 0),
		(drawing, 1334, 20, 2048, 30, 0),
		(drawing, 1335, 20, 2048, 30, 0),
		(drawing, 1336, 20, 2048, 30, 0),
		(drawing, 1337, 20, 2048, 30, 0),
		(drawing, 1338, 20, 2048, 30, 0),
		(drawing, 1339, 20, 2048, 30, 0),
		(drawing, 1340, 20, 2048, 30, 0),
		(drawing, 1341, 20, 2048, 30, 0),
		(drawing, 1342, 20, 2048, 30, 0),
		(drawing, 1343, 20, 2048, 30, 0),
		(drawing, 1344, 20, 2048, 30, 0),
		(drawing, 1345, 20, 2048, 30, 0),
		(drawing, 1346, 20, 2048, 30, 0),
		(drawing, 1347, 20, 2048, 30, 0),
		(drawing, 1348, 20, 2048, 30, 0),
		(drawing, 1349, 20, 2048, 30, 0),
		(drawing, 1350, 20, 2048, 30, 0),
		(drawing, 1351, 20, 2048, 30, 0),
		(drawing, 1352, 20, 2048, 30, 0),
		(drawing, 1353, 20, 2048, 30, 0),
		(drawing, 1354, 20, 2048, 30, 0),
		(drawing, 1355, 20, 2048, 30, 0),
		(drawing, 1356, 20, 2048, 30, 0),
		(drawing, 1357, 20, 2048, 30, 0),
		(drawing, 1358, 20, 2048, 30, 0),
		(drawing, 1359, 20, 2048, 30, 0),
		(drawing, 1360, 20, 2048, 30, 0),
		(drawing, 1361, 20, 2048, 30, 0),
		(drawing, 1362, 20, 2048, 30, 0),
		(drawing, 1363, 20, 2048, 30, 0),
		(drawing, 1364, 20, 2048, 30, 0),
		(drawing, 1365, 20, 2048, 30, 0),
		(drawing, 1366, 20, 2048, 30, 0),
		(drawing, 1367, 20, 2048, 30, 0),
		(drawing, 1368, 20, 2048, 30, 0),
		(drawing, 1369, 20, 2048, 30, 0),
		(drawing, 1370, 20, 2048, 30, 0),
		(drawing, 1371, 20, 2048, 30, 0),
		(drawing, 1372, 20, 2048, 30, 0),
		(drawing, 1373, 20, 2048, 30, 0),
		(drawing, 1374, 20, 2048, 30, 0),
		(drawing, 1375, 20, 2048, 30, 0),
		(drawing, 1376, 20, 2048, 30, 0),
		(drawing, 1377, 20, 2048, 30, 0),
		(drawing, 1378, 20, 2048, 30, 0),
		(drawing, 1379, 20, 2048, 30, 0),
		(drawing, 1380, 20, 2048, 30, 0),
		(drawing, 1381, 20, 2048, 30, 0),
		(drawing, 1382, 20, 2048, 30, 0),
		(drawing, 1383, 20, 2048, 30, 0),
		(drawing, 1384, 20, 2048, 30, 0),
		(drawing, 1385, 20, 2048, 30, 0),
		(drawing, 1386, 20, 2048, 30, 0),
		(drawing, 1387, 20, 2048, 30, 0),
		(drawing, 1388, 20, 2048, 30, 0),
		(drawing, 1389, 20, 2048, 30, 0),
		(drawing, 1390, 20, 2048, 30, 0),
		(drawing, 1391, 20, 2048, 30, 0),
		(drawing, 1392, 20, 2048, 30, 0),
		(drawing, 1393, 20, 2048, 30, 0),
		(drawing, 1394, 20, 2048, 30, 0),
		(drawing, 1395, 20, 2048, 30, 0),
		(drawing, 1396, 20, 2048, 30, 0),
		(drawing, 1397, 20, 2048, 30, 0),
		(drawing, 1398, 20, 2048, 30, 0),
		(drawing, 1399, 20, 2048, 30, 0),
		(drawing, 1400, 21, 2048, 30, 0),
		(drawing, 1401, 21, 2048, 30, 0),
		(drawing, 1402, 21, 2048, 30, 0),
		(drawing, 1403, 21, 2048, 30, 0),
		(drawing, 1404, 21, 2048, 30, 0),
		(drawing, 1405, 21, 2048, 30, 0),
		(drawing, 1406, 21, 2048, 30, 0),
		(drawing, 1407, 21, 2048, 30, 0),
		(drawing, 1408, 21, 2048, 30, 0),
		(drawing, 1409, 21, 2048, 30, 0),
		(drawing, 1410, 21, 2048, 30, 0),
		(drawing, 1411, 21, 2048, 30, 0),
		(drawing, 1412, 21, 2048, 30, 0),
		(drawing, 1413, 21, 2048, 30, 0),
		(drawing, 1414, 21, 2048, 30, 0),
		(drawing, 1415, 21, 2048, 30, 0),
		(drawing, 1416, 21, 2048, 30, 0),
		(drawing, 1417, 21, 2048, 30, 0),
		(drawing, 1418, 21, 2048, 30, 0),
		(drawing, 1419, 21, 2048, 30, 0),
		(drawing, 1420, 21, 2048, 30, 0),
		(drawing, 1421, 21, 2048, 30, 0),
		(drawing, 1422, 21, 2048, 30, 0),
		(drawing, 1423, 21, 2048, 30, 0),
		(drawing, 1424, 21, 2048, 30, 0),
		(drawing, 1425, 21, 2048, 30, 0),
		(drawing, 1426, 21, 2048, 30, 0),
		(drawing, 1427, 21, 2048, 30, 0),
		(drawing, 1428, 21, 2048, 30, 0),
		(drawing, 1429, 21, 2048, 30, 0),
		(drawing, 1430, 21, 2048, 30, 0),
		(drawing, 1431, 21, 2048, 30, 0),
		(drawing, 1432, 21, 2048, 30, 0),
		(drawing, 1433, 21, 2048, 30, 0),
		(drawing, 1434, 21, 2048, 30, 0),
		(drawing, 1435, 21, 2048, 30, 0),
		(drawing, 1436, 21, 2048, 30, 0),
		(drawing, 1437, 21, 2048, 30, 0),
		(drawing, 1438, 21, 2048, 30, 0),
		(drawing, 1439, 21, 2048, 30, 0),
		(drawing, 1440, 21, 2048, 30, 0),
		(drawing, 1441, 21, 2048, 30, 0),
		(drawing, 1442, 21, 2048, 30, 0),
		(drawing, 1443, 21, 2048, 30, 0),
		(drawing, 1444, 21, 2048, 30, 0),
		(drawing, 1445, 21, 2048, 30, 0),
		(drawing, 1446, 21, 2048, 30, 0),
		(drawing, 1447, 21, 2048, 30, 0),
		(drawing, 1448, 21, 2048, 30, 0),
		(drawing, 1449, 21, 2048, 30, 0),
		(drawing, 1450, 21, 2048, 30, 0),
		(drawing, 1451, 21, 2048, 30, 0),
		(drawing, 1452, 21, 2048, 30, 0),
		(drawing, 1453, 21, 2048, 30, 0),
		(drawing, 1454, 21, 2048, 30, 0),
		(drawing, 1455, 21, 2048, 30, 0),
		(drawing, 1456, 21, 2048, 30, 0),
		(drawing, 1457, 21, 2048, 30, 0),
		(drawing, 1458, 21, 2048, 30, 0),
		(drawing, 1459, 21, 2048, 30, 0),
		(drawing, 1460, 21, 2048, 30, 0),
		(drawing, 1461, 21, 2048, 30, 0),
		(drawing, 1462, 21, 2048, 30, 0),
		(drawing, 1463, 21, 2048, 30, 0),
		(drawing, 1464, 21, 2048, 30, 0),
		(drawing, 1465, 21, 2048, 30, 0),
		(drawing, 1466, 21, 2048, 30, 0),
		(drawing, 1467, 21, 2048, 30, 0),
		(drawing, 1468, 22, 2048, 30, 0),
		(drawing, 1469, 22, 2048, 30, 0),
		(drawing, 1470, 22, 2048, 30, 0),
		(drawing, 1471, 22, 2048, 30, 0),
		(drawing, 1472, 22, 2048, 30, 0),
		(drawing, 1473, 22, 2048, 30, 0),
		(drawing, 1474, 22, 2048, 30, 0),
		(drawing, 1475, 22, 2048, 30, 0),
		(drawing, 1476, 22, 2048, 30, 0),
		(drawing, 1477, 22, 2048, 30, 0),
		(drawing, 1478, 22, 2048, 30, 0),
		(drawing, 1479, 22, 2048, 30, 0),
		(drawing, 1480, 22, 2048, 30, 0),
		(drawing, 1481, 22, 2048, 30, 0),
		(drawing, 1482, 22, 2048, 30, 0),
		(drawing, 1483, 22, 2048, 30, 0),
		(drawing, 1484, 22, 2048, 30, 0),
		(drawing, 1485, 22, 2048, 30, 0),
		(drawing, 1486, 22, 2048, 30, 0),
		(drawing, 1487, 22, 2048, 30, 0),
		(drawing, 1488, 22, 2048, 30, 0),
		(drawing, 1489, 22, 2048, 30, 0),
		(drawing, 1490, 22, 2048, 30, 0),
		(drawing, 1491, 22, 2048, 30, 0),
		(drawing, 1492, 22, 2048, 30, 0),
		(drawing, 1493, 22, 2048, 30, 0),
		(drawing, 1494, 22, 2048, 30, 0),
		(drawing, 1495, 22, 2048, 30, 0),
		(drawing, 1496, 22, 2048, 30, 0),
		(drawing, 1497, 22, 2048, 30, 0),
		(drawing, 1498, 22, 2048, 30, 0),
		(drawing, 1499, 22, 2048, 30, 0),
		(drawing, 1500, 22, 2048, 30, 0),
		(drawing, 1501, 22, 2048, 30, 0),
		(drawing, 1502, 22, 2048, 30, 0),
		(drawing, 1503, 22, 2048, 30, 0),
		(drawing, 1504, 22, 2048, 30, 0),
		(drawing, 1505, 22, 2048, 30, 0),
		(drawing, 1506, 22, 2048, 30, 0),
		(drawing, 1507, 22, 2048, 30, 0),
		(drawing, 1508, 22, 2048, 30, 0),
		(drawing, 1509, 22, 2048, 30, 0),
		(drawing, 1510, 22, 2048, 30, 0),
		(drawing, 1511, 22, 2048, 30, 0),
		(drawing, 1512, 22, 2048, 30, 0),
		(drawing, 1513, 22, 2048, 30, 0),
		(drawing, 1514, 22, 2048, 30, 0),
		(drawing, 1515, 22, 2048, 30, 0),
		(drawing, 1516, 22, 2048, 30, 0),
		(drawing, 1517, 22, 2048, 30, 0),
		(drawing, 1518, 22, 2048, 30, 0),
		(drawing, 1519, 22, 2048, 30, 0),
		(drawing, 1520, 22, 2048, 30, 0),
		(drawing, 1521, 22, 2048, 30, 0),
		(drawing, 1522, 22, 2048, 30, 0),
		(drawing, 1523, 22, 2048, 30, 0),
		(drawing, 1524, 22, 2048, 30, 0),
		(drawing, 1525, 22, 2048, 30, 0),
		(drawing, 1526, 22, 2048, 30, 0),
		(drawing, 1527, 22, 2048, 30, 0),
		(drawing, 1528, 22, 2048, 30, 0),
		(drawing, 1529, 22, 2048, 30, 0),
		(drawing, 1530, 22, 2048, 30, 0),
		(drawing, 1531, 22, 2048, 30, 0),
		(drawing, 1532, 22, 2048, 30, 0),
		(drawing, 1533, 22, 2048, 30, 0),
		(drawing, 1534, 22, 2048, 30, 0),
		(drawing, 1535, 22, 2048, 30, 0),
		(drawing, 1536, 23, 2048, 30, 0),
		(drawing, 1537, 23, 2048, 30, 0),
		(drawing, 1538, 23, 2048, 30, 0),
		(drawing, 1539, 23, 2048, 30, 0),
		(drawing, 1540, 23, 2048, 30, 0),
		(drawing, 1541, 23, 2048, 30, 0),
		(drawing, 1542, 23, 2048, 30, 0),
		(drawing, 1543, 23, 2048, 30, 0),
		(drawing, 1544, 23, 2048, 30, 0),
		(drawing, 1545, 23, 2048, 30, 0),
		(drawing, 1546, 23, 2048, 30, 0),
		(drawing, 1547, 23, 2048, 30, 0),
		(drawing, 1548, 23, 2048, 30, 0),
		(drawing, 1549, 23, 2048, 30, 0),
		(drawing, 1550, 23, 2048, 30, 0),
		(drawing, 1551, 23, 2048, 30, 0),
		(drawing, 1552, 23, 2048, 30, 0),
		(drawing, 1553, 23, 2048, 30, 0),
		(drawing, 1554, 23, 2048, 30, 0),
		(drawing, 1555, 23, 2048, 30, 0),
		(drawing, 1556, 23, 2048, 30, 0),
		(drawing, 1557, 23, 2048, 30, 0),
		(drawing, 1558, 23, 2048, 30, 0),
		(drawing, 1559, 23, 2048, 30, 0),
		(drawing, 1560, 23, 2048, 30, 0),
		(drawing, 1561, 23, 2048, 30, 0),
		(drawing, 1562, 23, 2048, 30, 0),
		(drawing, 1563, 23, 2048, 30, 0),
		(drawing, 1564, 23, 2048, 30, 0),
		(drawing, 1565, 23, 2048, 30, 0),
		(drawing, 1566, 23, 2048, 30, 0),
		(drawing, 1567, 23, 2048, 30, 0),
		(drawing, 1568, 23, 2048, 30, 0),
		(drawing, 1569, 23, 2048, 30, 0),
		(drawing, 1570, 23, 2048, 30, 0),
		(drawing, 1571, 23, 2048, 30, 0),
		(drawing, 1572, 23, 2048, 30, 0),
		(drawing, 1573, 23, 2048, 30, 0),
		(drawing, 1574, 23, 2048, 30, 0),
		(drawing, 1575, 23, 2048, 30, 0),
		(drawing, 1576, 23, 2048, 30, 0),
		(drawing, 1577, 23, 2048, 30, 0),
		(drawing, 1578, 23, 2048, 30, 0),
		(drawing, 1579, 23, 2048, 30, 0),
		(drawing, 1580, 23, 2048, 30, 0),
		(drawing, 1581, 23, 2048, 30, 0),
		(drawing, 1582, 23, 2048, 30, 0),
		(drawing, 1583, 23, 2048, 30, 0),
		(drawing, 1584, 23, 2048, 30, 0),
		(drawing, 1585, 23, 2048, 30, 0),
		(drawing, 1586, 23, 2048, 30, 0),
		(drawing, 1587, 23, 2048, 30, 0),
		(drawing, 1588, 23, 2048, 30, 0),
		(drawing, 1589, 23, 2048, 30, 0),
		(drawing, 1590, 23, 2048, 30, 0),
		(drawing, 1591, 23, 2048, 30, 0),
		(drawing, 1592, 23, 2048, 30, 0),
		(drawing, 1593, 23, 2048, 30, 0),
		(drawing, 1594, 23, 2048, 30, 0),
		(drawing, 1595, 23, 2048, 30, 0),
		(drawing, 1596, 23, 2048, 30, 0),
		(drawing, 1597, 23, 2048, 30, 0),
		(drawing, 1598, 23, 2048, 30, 0),
		(drawing, 1599, 23, 2048, 30, 0),
		(drawing, 1600, 23, 2048, 30, 0),
		(drawing, 1601, 23, 2048, 30, 0),
		(drawing, 1602, 23, 2048, 30, 0),
		(drawing, 1603, 23, 2048, 30, 0),
		(drawing, 1604, 23, 2048, 30, 0),
		(drawing, 1605, 24, 2048, 30, 0),
		(drawing, 1606, 24, 2048, 30, 0),
		(drawing, 1607, 24, 2048, 30, 0),
		(drawing, 1608, 24, 2048, 30, 0),
		(drawing, 1609, 24, 2048, 30, 0),
		(drawing, 1610, 24, 2048, 30, 0),
		(drawing, 1611, 24, 2048, 30, 0),
		(drawing, 1612, 24, 2048, 30, 0),
		(drawing, 1613, 24, 2048, 30, 0),
		(drawing, 1614, 24, 2048, 30, 0),
		(drawing, 1615, 24, 2048, 30, 0),
		(drawing, 1616, 24, 2048, 30, 0),
		(drawing, 1617, 24, 2048, 30, 0),
		(drawing, 1618, 24, 2048, 30, 0),
		(drawing, 1619, 24, 2048, 30, 0),
		(drawing, 1620, 24, 2048, 30, 0),
		(drawing, 1621, 24, 2048, 30, 0),
		(drawing, 1622, 24, 2048, 30, 0),
		(drawing, 1623, 24, 2048, 30, 0),
		(drawing, 1624, 24, 2048, 30, 0),
		(drawing, 1625, 24, 2048, 30, 0),
		(drawing, 1626, 24, 2048, 30, 0),
		(drawing, 1627, 24, 2048, 30, 0),
		(drawing, 1628, 24, 2048, 30, 0),
		(drawing, 1629, 24, 2048, 30, 0),
		(drawing, 1630, 24, 2048, 30, 0),
		(drawing, 1631, 24, 2048, 30, 0),
		(drawing, 1632, 24, 2048, 30, 0),
		(drawing, 1633, 24, 2048, 30, 0),
		(drawing, 1634, 24, 2048, 30, 0),
		(drawing, 1635, 24, 2048, 30, 0),
		(drawing, 1636, 24, 2048, 30, 0),
		(drawing, 1637, 24, 2048, 30, 0),
		(drawing, 1638, 24, 2048, 30, 0),
		(drawing, 1639, 24, 2048, 30, 0),
		(drawing, 1640, 24, 2048, 30, 0),
		(drawing, 1641, 24, 2048, 30, 0),
		(drawing, 1642, 24, 2048, 30, 0),
		(drawing, 1643, 24, 2048, 30, 0),
		(drawing, 1644, 24, 2048, 30, 0),
		(drawing, 1645, 24, 2048, 30, 0),
		(drawing, 1646, 24, 2048, 30, 0),
		(drawing, 1647, 24, 2048, 30, 0),
		(drawing, 1648, 24, 2048, 30, 0),
		(drawing, 1649, 24, 2048, 30, 0),
		(drawing, 1650, 24, 2048, 30, 0),
		(drawing, 1651, 24, 2048, 30, 0),
		(drawing, 1652, 24, 2048, 30, 0),
		(drawing, 1653, 24, 2048, 30, 0),
		(drawing, 1654, 24, 2048, 30, 0),
		(drawing, 1655, 24, 2048, 30, 0),
		(drawing, 1656, 24, 2048, 30, 0),
		(drawing, 1657, 24, 2048, 30, 0),
		(drawing, 1658, 24, 2048, 30, 0),
		(drawing, 1659, 24, 2048, 30, 0),
		(drawing, 1660, 24, 2048, 30, 0),
		(drawing, 1661, 24, 2048, 30, 0),
		(drawing, 1662, 24, 2048, 30, 0),
		(drawing, 1663, 24, 2048, 30, 0),
		(drawing, 1664, 24, 2048, 30, 0),
		(drawing, 1665, 24, 2048, 30, 0),
		(drawing, 1666, 24, 2048, 30, 0),
		(drawing, 1667, 24, 2048, 30, 0),
		(drawing, 1668, 24, 2048, 30, 0),
		(drawing, 1669, 24, 2048, 30, 0),
		(drawing, 1670, 24, 2048, 30, 0),
		(drawing, 1671, 24, 2048, 30, 0),
		(drawing, 1672, 24, 2048, 30, 0),
		(drawing, 1673, 25, 2048, 30, 0),
		(drawing, 1674, 25, 2048, 30, 0),
		(drawing, 1675, 25, 2048, 30, 0),
		(drawing, 1676, 25, 2048, 30, 0),
		(drawing, 1677, 25, 2048, 30, 0),
		(drawing, 1678, 25, 2048, 30, 0),
		(drawing, 1679, 25, 2048, 30, 0),
		(drawing, 1680, 25, 2048, 30, 0),
		(drawing, 1681, 25, 2048, 30, 0),
		(drawing, 1682, 25, 2048, 30, 0),
		(drawing, 1683, 25, 2048, 30, 0),
		(drawing, 1684, 25, 2048, 30, 0),
		(drawing, 1685, 25, 2048, 30, 0),
		(drawing, 1686, 25, 2048, 30, 0),
		(drawing, 1687, 25, 2048, 30, 0),
		(drawing, 1688, 25, 2048, 30, 0),
		(drawing, 1689, 25, 2048, 30, 0),
		(drawing, 1690, 25, 2048, 30, 0),
		(drawing, 1691, 25, 2048, 30, 0),
		(drawing, 1692, 25, 2048, 30, 0),
		(drawing, 1693, 25, 2048, 30, 0),
		(drawing, 1694, 25, 2048, 30, 0),
		(drawing, 1695, 25, 2048, 30, 0),
		(drawing, 1696, 25, 2048, 30, 0),
		(drawing, 1697, 25, 2048, 30, 0),
		(drawing, 1698, 25, 2048, 30, 0),
		(drawing, 1699, 25, 2048, 30, 0),
		(drawing, 1700, 25, 2048, 30, 0),
		(drawing, 1701, 25, 2048, 30, 0),
		(drawing, 1702, 25, 2048, 30, 0),
		(drawing, 1703, 25, 2048, 30, 0),
		(drawing, 1704, 25, 2048, 30, 0),
		(drawing, 1705, 25, 2048, 30, 0),
		(drawing, 1706, 25, 2048, 30, 0),
		(drawing, 1707, 25, 2048, 30, 0),
		(drawing, 1708, 25, 2048, 30, 0),
		(drawing, 1709, 25, 2048, 30, 0),
		(drawing, 1710, 25, 2048, 30, 0),
		(drawing, 1711, 25, 2048, 30, 0),
		(drawing, 1712, 25, 2048, 30, 0),
		(drawing, 1713, 25, 2048, 30, 0),
		(drawing, 1714, 25, 2048, 30, 0),
		(drawing, 1715, 25, 2048, 30, 0),
		(drawing, 1716, 25, 2048, 30, 0),
		(drawing, 1717, 25, 2048, 30, 0),
		(drawing, 1718, 25, 2048, 30, 0),
		(drawing, 1719, 25, 2048, 30, 0),
		(drawing, 1720, 25, 2048, 30, 0),
		(drawing, 1721, 25, 2048, 30, 0),
		(drawing, 1722, 25, 2048, 30, 0),
		(drawing, 1723, 25, 2048, 30, 0),
		(drawing, 1724, 25, 2048, 30, 0),
		(drawing, 1725, 25, 2048, 30, 0),
		(drawing, 1726, 25, 2048, 30, 0),
		(drawing, 1727, 25, 2048, 30, 0),
		(drawing, 1728, 25, 2048, 30, 0),
		(drawing, 1729, 25, 2048, 30, 0),
		(drawing, 1730, 25, 2048, 30, 0),
		(drawing, 1731, 25, 2048, 30, 0),
		(drawing, 1732, 25, 2048, 30, 0),
		(drawing, 1733, 25, 2048, 30, 0),
		(drawing, 1734, 25, 2048, 30, 0),
		(drawing, 1735, 25, 2048, 30, 0),
		(drawing, 1736, 25, 2048, 30, 0),
		(drawing, 1737, 25, 2048, 30, 0),
		(drawing, 1738, 25, 2048, 30, 0),
		(drawing, 1739, 25, 2048, 30, 0),
		(drawing, 1740, 25, 2048, 30, 0),
		(drawing, 1741, 26, 2048, 30, 0),
		(drawing, 1742, 26, 2048, 30, 0),
		(drawing, 1743, 26, 2048, 30, 0),
		(drawing, 1744, 26, 2048, 30, 0),
		(drawing, 1745, 26, 2048, 30, 0),
		(drawing, 1746, 26, 2048, 30, 0),
		(drawing, 1747, 26, 2048, 30, 0),
		(drawing, 1748, 26, 2048, 30, 0),
		(drawing, 1749, 26, 2048, 30, 0),
		(drawing, 1750, 26, 2048, 30, 0),
		(drawing, 1751, 26, 2048, 30, 0),
		(drawing, 1752, 26, 2048, 30, 0),
		(drawing, 1753, 26, 2048, 30, 0),
		(drawing, 1754, 26, 2048, 30, 0),
		(drawing, 1755, 26, 2048, 30, 0),
		(drawing, 1756, 26, 2048, 30, 0),
		(drawing, 1757, 26, 2048, 30, 0),
		(drawing, 1758, 26, 2048, 30, 0),
		(drawing, 1759, 26, 2048, 30, 0),
		(drawing, 1760, 26, 2048, 30, 0),
		(drawing, 1761, 26, 2048, 30, 0),
		(drawing, 1762, 26, 2048, 30, 0),
		(drawing, 1763, 26, 2048, 30, 0),
		(drawing, 1764, 26, 2048, 30, 0),
		(drawing, 1765, 26, 2048, 30, 0),
		(drawing, 1766, 26, 2048, 30, 0),
		(drawing, 1767, 26, 2048, 30, 0),
		(drawing, 1768, 26, 2048, 30, 0),
		(drawing, 1769, 26, 2048, 30, 0),
		(drawing, 1770, 26, 2048, 30, 0),
		(drawing, 1771, 26, 2048, 30, 0),
		(drawing, 1772, 26, 2048, 30, 0),
		(drawing, 1773, 26, 2048, 30, 0),
		(drawing, 1774, 26, 2048, 30, 0),
		(drawing, 1775, 26, 2048, 30, 0),
		(drawing, 1776, 26, 2048, 30, 0),
		(drawing, 1777, 26, 2048, 30, 0),
		(drawing, 1778, 26, 2048, 30, 0),
		(drawing, 1779, 26, 2048, 30, 0),
		(drawing, 1780, 26, 2048, 30, 0),
		(drawing, 1781, 26, 2048, 30, 0),
		(drawing, 1782, 26, 2048, 30, 0),
		(drawing, 1783, 26, 2048, 30, 0),
		(drawing, 1784, 26, 2048, 30, 0),
		(drawing, 1785, 26, 2048, 30, 0),
		(drawing, 1786, 26, 2048, 30, 0),
		(drawing, 1787, 26, 2048, 30, 0),
		(drawing, 1788, 26, 2048, 30, 0),
		(drawing, 1789, 26, 2048, 30, 0),
		(drawing, 1790, 26, 2048, 30, 0),
		(drawing, 1791, 26, 2048, 30, 0),
		(drawing, 1792, 26, 2048, 30, 0),
		(drawing, 1793, 26, 2048, 30, 0),
		(drawing, 1794, 26, 2048, 30, 0),
		(drawing, 1795, 26, 2048, 30, 0),
		(drawing, 1796, 26, 2048, 30, 0),
		(drawing, 1797, 26, 2048, 30, 0),
		(drawing, 1798, 26, 2048, 30, 0),
		(drawing, 1799, 26, 2048, 30, 0),
		(drawing, 1800, 26, 2048, 30, 0),
		(drawing, 1801, 26, 2048, 30, 0),
		(drawing, 1802, 26, 2048, 30, 0),
		(drawing, 1803, 26, 2048, 30, 0),
		(drawing, 1804, 26, 2048, 30, 0),
		(drawing, 1805, 26, 2048, 30, 0),
		(drawing, 1806, 26, 2048, 30, 0),
		(drawing, 1807, 26, 2048, 30, 0),
		(drawing, 1808, 26, 2048, 30, 0),
		(drawing, 1809, 26, 2048, 30, 0),
		(drawing, 1810, 27, 2048, 30, 0),
		(drawing, 1811, 27, 2048, 30, 0),
		(drawing, 1812, 27, 2048, 30, 0),
		(drawing, 1813, 27, 2048, 30, 0),
		(drawing, 1814, 27, 2048, 30, 0),
		(drawing, 1815, 27, 2048, 30, 0),
		(drawing, 1816, 27, 2048, 30, 0),
		(drawing, 1817, 27, 2048, 30, 0),
		(drawing, 1818, 27, 2048, 30, 0),
		(drawing, 1819, 27, 2048, 30, 0),
		(drawing, 1820, 27, 2048, 30, 0),
		(drawing, 1821, 27, 2048, 30, 0),
		(drawing, 1822, 27, 2048, 30, 0),
		(drawing, 1823, 27, 2048, 30, 0),
		(drawing, 1824, 27, 2048, 30, 0),
		(drawing, 1825, 27, 2048, 30, 0),
		(drawing, 1826, 27, 2048, 30, 0),
		(drawing, 1827, 27, 2048, 30, 0),
		(drawing, 1828, 27, 2048, 30, 0),
		(drawing, 1829, 27, 2048, 30, 0),
		(drawing, 1830, 27, 2048, 30, 0),
		(drawing, 1831, 27, 2048, 30, 0),
		(drawing, 1832, 27, 2048, 30, 0),
		(drawing, 1833, 27, 2048, 30, 0),
		(drawing, 1834, 27, 2048, 30, 0),
		(drawing, 1835, 27, 2048, 30, 0),
		(drawing, 1836, 27, 2048, 30, 0),
		(drawing, 1837, 27, 2048, 30, 0),
		(drawing, 1838, 27, 2048, 30, 0),
		(drawing, 1839, 27, 2048, 30, 0),
		(drawing, 1840, 27, 2048, 30, 0),
		(drawing, 1841, 27, 2048, 30, 0),
		(drawing, 1842, 27, 2048, 30, 0),
		(drawing, 1843, 27, 2048, 30, 0),
		(drawing, 1844, 27, 2048, 30, 0),
		(drawing, 1845, 27, 2048, 30, 0),
		(drawing, 1846, 27, 2048, 30, 0),
		(drawing, 1847, 27, 2048, 30, 0),
		(drawing, 1848, 27, 2048, 30, 0),
		(drawing, 1849, 27, 2048, 30, 0),
		(drawing, 1850, 27, 2048, 30, 0),
		(drawing, 1851, 27, 2048, 30, 0),
		(drawing, 1852, 27, 2048, 30, 0),
		(drawing, 1853, 27, 2048, 30, 0),
		(drawing, 1854, 27, 2048, 30, 0),
		(drawing, 1855, 27, 2048, 30, 0),
		(drawing, 1856, 27, 2048, 30, 0),
		(drawing, 1857, 27, 2048, 30, 0),
		(drawing, 1858, 27, 2048, 30, 0),
		(drawing, 1859, 27, 2048, 30, 0),
		(drawing, 1860, 27, 2048, 30, 0),
		(drawing, 1861, 27, 2048, 30, 0),
		(drawing, 1862, 27, 2048, 30, 0),
		(drawing, 1863, 27, 2048, 30, 0),
		(drawing, 1864, 27, 2048, 30, 0),
		(drawing, 1865, 27, 2048, 30, 0),
		(drawing, 1866, 27, 2048, 30, 0),
		(drawing, 1867, 27, 2048, 30, 0),
		(drawing, 1868, 27, 2048, 30, 0),
		(drawing, 1869, 27, 2048, 30, 0),
		(drawing, 1870, 27, 2048, 30, 0),
		(drawing, 1871, 27, 2048, 30, 0),
		(drawing, 1872, 27, 2048, 30, 0),
		(drawing, 1873, 27, 2048, 30, 0),
		(drawing, 1874, 27, 2048, 30, 0),
		(drawing, 1875, 27, 2048, 30, 0),
		(drawing, 1876, 27, 2048, 30, 0),
		(drawing, 1877, 27, 2048, 30, 0),
		(drawing, 1878, 28, 2048, 30, 0),
		(drawing, 1879, 28, 2048, 30, 0),
		(drawing, 1880, 28, 2048, 30, 0),
		(drawing, 1881, 28, 2048, 30, 0),
		(drawing, 1882, 28, 2048, 30, 0),
		(drawing, 1883, 28, 2048, 30, 0),
		(drawing, 1884, 28, 2048, 30, 0),
		(drawing, 1885, 28, 2048, 30, 0),
		(drawing, 1886, 28, 2048, 30, 0),
		(drawing, 1887, 28, 2048, 30, 0),
		(drawing, 1888, 28, 2048, 30, 0),
		(drawing, 1889, 28, 2048, 30, 0),
		(drawing, 1890, 28, 2048, 30, 0),
		(drawing, 1891, 28, 2048, 30, 0),
		(drawing, 1892, 28, 2048, 30, 0),
		(drawing, 1893, 28, 2048, 30, 0),
		(drawing, 1894, 28, 2048, 30, 0),
		(drawing, 1895, 28, 2048, 30, 0),
		(drawing, 1896, 28, 2048, 30, 0),
		(drawing, 1897, 28, 2048, 30, 0),
		(drawing, 1898, 28, 2048, 30, 0),
		(drawing, 1899, 28, 2048, 30, 0),
		(drawing, 1900, 28, 2048, 30, 0),
		(drawing, 1901, 28, 2048, 30, 0),
		(drawing, 1902, 28, 2048, 30, 0),
		(drawing, 1903, 28, 2048, 30, 0),
		(drawing, 1904, 28, 2048, 30, 0),
		(drawing, 1905, 28, 2048, 30, 0),
		(drawing, 1906, 28, 2048, 30, 0),
		(drawing, 1907, 28, 2048, 30, 0),
		(drawing, 1908, 28, 2048, 30, 0),
		(drawing, 1909, 28, 2048, 30, 0),
		(drawing, 1910, 28, 2048, 30, 0),
		(drawing, 1911, 28, 2048, 30, 0),
		(drawing, 1912, 28, 2048, 30, 0),
		(drawing, 1913, 28, 2048, 30, 0),
		(drawing, 1914, 28, 2048, 30, 0),
		(drawing, 1915, 28, 2048, 30, 0),
		(drawing, 1916, 28, 2048, 30, 0),
		(drawing, 1917, 28, 2048, 30, 0),
		(drawing, 1918, 28, 2048, 30, 0),
		(drawing, 1919, 28, 2048, 30, 0),
		(drawing, 1920, 28, 2048, 30, 0),
		(drawing, 1921, 28, 2048, 30, 0),
		(drawing, 1922, 28, 2048, 30, 0),
		(drawing, 1923, 28, 2048, 30, 0),
		(drawing, 1924, 28, 2048, 30, 0),
		(drawing, 1925, 28, 2048, 30, 0),
		(drawing, 1926, 28, 2048, 30, 0),
		(drawing, 1927, 28, 2048, 30, 0),
		(drawing, 1928, 28, 2048, 30, 0),
		(drawing, 1929, 28, 2048, 30, 0),
		(drawing, 1930, 28, 2048, 30, 0),
		(drawing, 1931, 28, 2048, 30, 0),
		(drawing, 1932, 28, 2048, 30, 0),
		(drawing, 1933, 28, 2048, 30, 0),
		(drawing, 1934, 28, 2048, 30, 0),
		(drawing, 1935, 28, 2048, 30, 0),
		(drawing, 1936, 28, 2048, 30, 0),
		(drawing, 1937, 28, 2048, 30, 0),
		(drawing, 1938, 28, 2048, 30, 0),
		(drawing, 1939, 28, 2048, 30, 0),
		(drawing, 1940, 28, 2048, 30, 0),
		(drawing, 1941, 28, 2048, 30, 0),
		(drawing, 1942, 28, 2048, 30, 0),
		(drawing, 1943, 28, 2048, 30, 0),
		(drawing, 1944, 28, 2048, 30, 0),
		(drawing, 1945, 28, 2048, 30, 0),
		(drawing, 1946, 29, 2048, 30, 0),
		(drawing, 1947, 29, 2048, 30, 0),
		(drawing, 1948, 29, 2048, 30, 0),
		(drawing, 1949, 29, 2048, 30, 0),
		(drawing, 1950, 29, 2048, 30, 0),
		(drawing, 1951, 29, 2048, 30, 0),
		(drawing, 1952, 29, 2048, 30, 0),
		(drawing, 1953, 29, 2048, 30, 0),
		(drawing, 1954, 29, 2048, 30, 0),
		(drawing, 1955, 29, 2048, 30, 0),
		(drawing, 1956, 29, 2048, 30, 0),
		(drawing, 1957, 29, 2048, 30, 0),
		(drawing, 1958, 29, 2048, 30, 0),
		(drawing, 1959, 29, 2048, 30, 0),
		(drawing, 1960, 29, 2048, 30, 0),
		(drawing, 1961, 29, 2048, 30, 0),
		(drawing, 1962, 29, 2048, 30, 0),
		(drawing, 1963, 29, 2048, 30, 0),
		(drawing, 1964, 29, 2048, 30, 0),
		(drawing, 1965, 29, 2048, 30, 0),
		(drawing, 1966, 29, 2048, 30, 0),
		(drawing, 1967, 29, 2048, 30, 0),
		(drawing, 1968, 29, 2048, 30, 0),
		(drawing, 1969, 29, 2048, 30, 0),
		(drawing, 1970, 29, 2048, 30, 0),
		(drawing, 1971, 29, 2048, 30, 0),
		(drawing, 1972, 29, 2048, 30, 0),
		(drawing, 1973, 29, 2048, 30, 0),
		(drawing, 1974, 29, 2048, 30, 0),
		(drawing, 1975, 29, 2048, 30, 0),
		(drawing, 1976, 29, 2048, 30, 0),
		(drawing, 1977, 29, 2048, 30, 0),
		(drawing, 1978, 29, 2048, 30, 0),
		(drawing, 1979, 29, 2048, 30, 0),
		(drawing, 1980, 29, 2048, 30, 0),
		(drawing, 1981, 29, 2048, 30, 0),
		(drawing, 1982, 29, 2048, 30, 0),
		(drawing, 1983, 29, 2048, 30, 0),
		(drawing, 1984, 29, 2048, 30, 0),
		(drawing, 1985, 29, 2048, 30, 0),
		(drawing, 1986, 29, 2048, 30, 0),
		(drawing, 1987, 29, 2048, 30, 0),
		(drawing, 1988, 29, 2048, 30, 0),
		(drawing, 1989, 29, 2048, 30, 0),
		(drawing, 1990, 29, 2048, 30, 0),
		(drawing, 1991, 29, 2048, 30, 0),
		(drawing, 1992, 29, 2048, 30, 0),
		(drawing, 1993, 29, 2048, 30, 0),
		(drawing, 1994, 29, 2048, 30, 0),
		(drawing, 1995, 29, 2048, 30, 0),
		(drawing, 1996, 29, 2048, 30, 0),
		(drawing, 1997, 29, 2048, 30, 0),
		(drawing, 1998, 29, 2048, 30, 0),
		(drawing, 1999, 29, 2048, 30, 0),
		(drawing, 2000, 29, 2048, 30, 0),
		(drawing, 2001, 29, 2048, 30, 0),
		(drawing, 2002, 29, 2048, 30, 0),
		(drawing, 2003, 29, 2048, 30, 0),
		(drawing, 2004, 29, 2048, 30, 0),
		(drawing, 2005, 29, 2048, 30, 0),
		(drawing, 2006, 29, 2048, 30, 0),
		(drawing, 2007, 29, 2048, 30, 0),
		(drawing, 2008, 29, 2048, 30, 0),
		(drawing, 2009, 29, 2048, 30, 0),
		(drawing, 2010, 29, 2048, 30, 0),
		(drawing, 2011, 29, 2048, 30, 0),
		(drawing, 2012, 29, 2048, 30, 0),
		(drawing, 2013, 29, 2048, 30, 0),
		(drawing, 2014, 30, 2048, 30, 0),
		(drawing, 2015, 30, 2048, 30, 0),
		(drawing, 2016, 30, 2048, 30, 0),
		(drawing, 2017, 30, 2048, 30, 0),
		(drawing, 2018, 30, 2048, 30, 0),
		(drawing, 2019, 30, 2048, 30, 0),
		(drawing, 2020, 30, 2048, 30, 0),
		(drawing, 2021, 30, 2048, 30, 0),
		(drawing, 2022, 30, 2048, 30, 0),
		(drawing, 2023, 30, 2048, 30, 0),
		(drawing, 2024, 30, 2048, 30, 0),
		(drawing, 2025, 30, 2048, 30, 0),
		(drawing, 2026, 30, 2048, 30, 0),
		(drawing, 2027, 30, 2048, 30, 0),
		(drawing, 2028, 30, 2048, 30, 0),
		(drawing, 2029, 30, 2048, 30, 0),
		(drawing, 2030, 30, 2048, 30, 0),
		(drawing, 2031, 30, 2048, 30, 0),
		(drawing, 2032, 30, 2048, 30, 0),
		(drawing, 2033, 30, 2048, 30, 0),
		(drawing, 2034, 30, 2048, 30, 0),
		(drawing, 2035, 30, 2048, 30, 0),
		(drawing, 2036, 30, 2048, 30, 0),
		(drawing, 2037, 30, 2048, 30, 0),
		(drawing, 2038, 30, 2048, 30, 0),
		(drawing, 2039, 30, 2048, 30, 0),
		(drawing, 2040, 30, 2048, 30, 0),
		(drawing, 2041, 30, 2048, 30, 0),
		(drawing, 2042, 30, 2048, 30, 0),
		(drawing, 2043, 30, 2048, 30, 0),
		(drawing, 2044, 30, 2048, 30, 0),
		(drawing, 2045, 30, 2048, 30, 0),
		(drawing, 2046, 30, 2048, 30, 0),
		(drawing, 2047, 30, 2048, 30, 0),
		(done, 2048, 30, 2048, 30, 0)
	);
END PACKAGE ex1_data_pak;
