-- advanced test 6
-- draw line from (0,0) to (2048,0)
-- NOTE * xin,yin are 12bits logic vectors
--------* 2048 in decimal is b1000,0000,0000
--------* this test is for xincr= b1000,0000,0000


PACKAGE ex1_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        txt: cyc; --see above definition
        x,y: INTEGER;   -- x,y are pixel coordinate outputs
        xin,yin: INTEGER; -- xn,yn are inputs xin, yin (0-4095)
        xbias: INTEGER; -- input xbias (1 or 0)
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(

		(reset, 0, 0, 0, 0, 0),
		(start, 0, 0, 2048, 0, 0),
		(drawing, 0, 0, 2048, 0, 0),
		(drawing, 1, 0, 2048, 0, 0),
		(drawing, 2, 0, 2048, 0, 0),
		(drawing, 3, 0, 2048, 0, 0),
		(drawing, 4, 0, 2048, 0, 0),
		(drawing, 5, 0, 2048, 0, 0),
		(drawing, 6, 0, 2048, 0, 0),
		(drawing, 7, 0, 2048, 0, 0),
		(drawing, 8, 0, 2048, 0, 0),
		(drawing, 9, 0, 2048, 0, 0),
		(drawing, 10, 0, 2048, 0, 0),
		(drawing, 11, 0, 2048, 0, 0),
		(drawing, 12, 0, 2048, 0, 0),
		(drawing, 13, 0, 2048, 0, 0),
		(drawing, 14, 0, 2048, 0, 0),
		(drawing, 15, 0, 2048, 0, 0),
		(drawing, 16, 0, 2048, 0, 0),
		(drawing, 17, 0, 2048, 0, 0),
		(drawing, 18, 0, 2048, 0, 0),
		(drawing, 19, 0, 2048, 0, 0),
		(drawing, 20, 0, 2048, 0, 0),
		(drawing, 21, 0, 2048, 0, 0),
		(drawing, 22, 0, 2048, 0, 0),
		(drawing, 23, 0, 2048, 0, 0),
		(drawing, 24, 0, 2048, 0, 0),
		(drawing, 25, 0, 2048, 0, 0),
		(drawing, 26, 0, 2048, 0, 0),
		(drawing, 27, 0, 2048, 0, 0),
		(drawing, 28, 0, 2048, 0, 0),
		(drawing, 29, 0, 2048, 0, 0),
		(drawing, 30, 0, 2048, 0, 0),
		(drawing, 31, 0, 2048, 0, 0),
		(drawing, 32, 0, 2048, 0, 0),
		(drawing, 33, 0, 2048, 0, 0),
		(drawing, 34, 0, 2048, 0, 0),
		(drawing, 35, 0, 2048, 0, 0),
		(drawing, 36, 0, 2048, 0, 0),
		(drawing, 37, 0, 2048, 0, 0),
		(drawing, 38, 0, 2048, 0, 0),
		(drawing, 39, 0, 2048, 0, 0),
		(drawing, 40, 0, 2048, 0, 0),
		(drawing, 41, 0, 2048, 0, 0),
		(drawing, 42, 0, 2048, 0, 0),
		(drawing, 43, 0, 2048, 0, 0),
		(drawing, 44, 0, 2048, 0, 0),
		(drawing, 45, 0, 2048, 0, 0),
		(drawing, 46, 0, 2048, 0, 0),
		(drawing, 47, 0, 2048, 0, 0),
		(drawing, 48, 0, 2048, 0, 0),
		(drawing, 49, 0, 2048, 0, 0),
		(drawing, 50, 0, 2048, 0, 0),
		(drawing, 51, 0, 2048, 0, 0),
		(drawing, 52, 0, 2048, 0, 0),
		(drawing, 53, 0, 2048, 0, 0),
		(drawing, 54, 0, 2048, 0, 0),
		(drawing, 55, 0, 2048, 0, 0),
		(drawing, 56, 0, 2048, 0, 0),
		(drawing, 57, 0, 2048, 0, 0),
		(drawing, 58, 0, 2048, 0, 0),
		(drawing, 59, 0, 2048, 0, 0),
		(drawing, 60, 0, 2048, 0, 0),
		(drawing, 61, 0, 2048, 0, 0),
		(drawing, 62, 0, 2048, 0, 0),
		(drawing, 63, 0, 2048, 0, 0),
		(drawing, 64, 0, 2048, 0, 0),
		(drawing, 65, 0, 2048, 0, 0),
		(drawing, 66, 0, 2048, 0, 0),
		(drawing, 67, 0, 2048, 0, 0),
		(drawing, 68, 0, 2048, 0, 0),
		(drawing, 69, 0, 2048, 0, 0),
		(drawing, 70, 0, 2048, 0, 0),
		(drawing, 71, 0, 2048, 0, 0),
		(drawing, 72, 0, 2048, 0, 0),
		(drawing, 73, 0, 2048, 0, 0),
		(drawing, 74, 0, 2048, 0, 0),
		(drawing, 75, 0, 2048, 0, 0),
		(drawing, 76, 0, 2048, 0, 0),
		(drawing, 77, 0, 2048, 0, 0),
		(drawing, 78, 0, 2048, 0, 0),
		(drawing, 79, 0, 2048, 0, 0),
		(drawing, 80, 0, 2048, 0, 0),
		(drawing, 81, 0, 2048, 0, 0),
		(drawing, 82, 0, 2048, 0, 0),
		(drawing, 83, 0, 2048, 0, 0),
		(drawing, 84, 0, 2048, 0, 0),
		(drawing, 85, 0, 2048, 0, 0),
		(drawing, 86, 0, 2048, 0, 0),
		(drawing, 87, 0, 2048, 0, 0),
		(drawing, 88, 0, 2048, 0, 0),
		(drawing, 89, 0, 2048, 0, 0),
		(drawing, 90, 0, 2048, 0, 0),
		(drawing, 91, 0, 2048, 0, 0),
		(drawing, 92, 0, 2048, 0, 0),
		(drawing, 93, 0, 2048, 0, 0),
		(drawing, 94, 0, 2048, 0, 0),
		(drawing, 95, 0, 2048, 0, 0),
		(drawing, 96, 0, 2048, 0, 0),
		(drawing, 97, 0, 2048, 0, 0),
		(drawing, 98, 0, 2048, 0, 0),
		(drawing, 99, 0, 2048, 0, 0),
		(drawing, 100, 0, 2048, 0, 0),
		(drawing, 101, 0, 2048, 0, 0),
		(drawing, 102, 0, 2048, 0, 0),
		(drawing, 103, 0, 2048, 0, 0),
		(drawing, 104, 0, 2048, 0, 0),
		(drawing, 105, 0, 2048, 0, 0),
		(drawing, 106, 0, 2048, 0, 0),
		(drawing, 107, 0, 2048, 0, 0),
		(drawing, 108, 0, 2048, 0, 0),
		(drawing, 109, 0, 2048, 0, 0),
		(drawing, 110, 0, 2048, 0, 0),
		(drawing, 111, 0, 2048, 0, 0),
		(drawing, 112, 0, 2048, 0, 0),
		(drawing, 113, 0, 2048, 0, 0),
		(drawing, 114, 0, 2048, 0, 0),
		(drawing, 115, 0, 2048, 0, 0),
		(drawing, 116, 0, 2048, 0, 0),
		(drawing, 117, 0, 2048, 0, 0),
		(drawing, 118, 0, 2048, 0, 0),
		(drawing, 119, 0, 2048, 0, 0),
		(drawing, 120, 0, 2048, 0, 0),
		(drawing, 121, 0, 2048, 0, 0),
		(drawing, 122, 0, 2048, 0, 0),
		(drawing, 123, 0, 2048, 0, 0),
		(drawing, 124, 0, 2048, 0, 0),
		(drawing, 125, 0, 2048, 0, 0),
		(drawing, 126, 0, 2048, 0, 0),
		(drawing, 127, 0, 2048, 0, 0),
		(drawing, 128, 0, 2048, 0, 0),
		(drawing, 129, 0, 2048, 0, 0),
		(drawing, 130, 0, 2048, 0, 0),
		(drawing, 131, 0, 2048, 0, 0),
		(drawing, 132, 0, 2048, 0, 0),
		(drawing, 133, 0, 2048, 0, 0),
		(drawing, 134, 0, 2048, 0, 0),
		(drawing, 135, 0, 2048, 0, 0),
		(drawing, 136, 0, 2048, 0, 0),
		(drawing, 137, 0, 2048, 0, 0),
		(drawing, 138, 0, 2048, 0, 0),
		(drawing, 139, 0, 2048, 0, 0),
		(drawing, 140, 0, 2048, 0, 0),
		(drawing, 141, 0, 2048, 0, 0),
		(drawing, 142, 0, 2048, 0, 0),
		(drawing, 143, 0, 2048, 0, 0),
		(drawing, 144, 0, 2048, 0, 0),
		(drawing, 145, 0, 2048, 0, 0),
		(drawing, 146, 0, 2048, 0, 0),
		(drawing, 147, 0, 2048, 0, 0),
		(drawing, 148, 0, 2048, 0, 0),
		(drawing, 149, 0, 2048, 0, 0),
		(drawing, 150, 0, 2048, 0, 0),
		(drawing, 151, 0, 2048, 0, 0),
		(drawing, 152, 0, 2048, 0, 0),
		(drawing, 153, 0, 2048, 0, 0),
		(drawing, 154, 0, 2048, 0, 0),
		(drawing, 155, 0, 2048, 0, 0),
		(drawing, 156, 0, 2048, 0, 0),
		(drawing, 157, 0, 2048, 0, 0),
		(drawing, 158, 0, 2048, 0, 0),
		(drawing, 159, 0, 2048, 0, 0),
		(drawing, 160, 0, 2048, 0, 0),
		(drawing, 161, 0, 2048, 0, 0),
		(drawing, 162, 0, 2048, 0, 0),
		(drawing, 163, 0, 2048, 0, 0),
		(drawing, 164, 0, 2048, 0, 0),
		(drawing, 165, 0, 2048, 0, 0),
		(drawing, 166, 0, 2048, 0, 0),
		(drawing, 167, 0, 2048, 0, 0),
		(drawing, 168, 0, 2048, 0, 0),
		(drawing, 169, 0, 2048, 0, 0),
		(drawing, 170, 0, 2048, 0, 0),
		(drawing, 171, 0, 2048, 0, 0),
		(drawing, 172, 0, 2048, 0, 0),
		(drawing, 173, 0, 2048, 0, 0),
		(drawing, 174, 0, 2048, 0, 0),
		(drawing, 175, 0, 2048, 0, 0),
		(drawing, 176, 0, 2048, 0, 0),
		(drawing, 177, 0, 2048, 0, 0),
		(drawing, 178, 0, 2048, 0, 0),
		(drawing, 179, 0, 2048, 0, 0),
		(drawing, 180, 0, 2048, 0, 0),
		(drawing, 181, 0, 2048, 0, 0),
		(drawing, 182, 0, 2048, 0, 0),
		(drawing, 183, 0, 2048, 0, 0),
		(drawing, 184, 0, 2048, 0, 0),
		(drawing, 185, 0, 2048, 0, 0),
		(drawing, 186, 0, 2048, 0, 0),
		(drawing, 187, 0, 2048, 0, 0),
		(drawing, 188, 0, 2048, 0, 0),
		(drawing, 189, 0, 2048, 0, 0),
		(drawing, 190, 0, 2048, 0, 0),
		(drawing, 191, 0, 2048, 0, 0),
		(drawing, 192, 0, 2048, 0, 0),
		(drawing, 193, 0, 2048, 0, 0),
		(drawing, 194, 0, 2048, 0, 0),
		(drawing, 195, 0, 2048, 0, 0),
		(drawing, 196, 0, 2048, 0, 0),
		(drawing, 197, 0, 2048, 0, 0),
		(drawing, 198, 0, 2048, 0, 0),
		(drawing, 199, 0, 2048, 0, 0),
		(drawing, 200, 0, 2048, 0, 0),
		(drawing, 201, 0, 2048, 0, 0),
		(drawing, 202, 0, 2048, 0, 0),
		(drawing, 203, 0, 2048, 0, 0),
		(drawing, 204, 0, 2048, 0, 0),
		(drawing, 205, 0, 2048, 0, 0),
		(drawing, 206, 0, 2048, 0, 0),
		(drawing, 207, 0, 2048, 0, 0),
		(drawing, 208, 0, 2048, 0, 0),
		(drawing, 209, 0, 2048, 0, 0),
		(drawing, 210, 0, 2048, 0, 0),
		(drawing, 211, 0, 2048, 0, 0),
		(drawing, 212, 0, 2048, 0, 0),
		(drawing, 213, 0, 2048, 0, 0),
		(drawing, 214, 0, 2048, 0, 0),
		(drawing, 215, 0, 2048, 0, 0),
		(drawing, 216, 0, 2048, 0, 0),
		(drawing, 217, 0, 2048, 0, 0),
		(drawing, 218, 0, 2048, 0, 0),
		(drawing, 219, 0, 2048, 0, 0),
		(drawing, 220, 0, 2048, 0, 0),
		(drawing, 221, 0, 2048, 0, 0),
		(drawing, 222, 0, 2048, 0, 0),
		(drawing, 223, 0, 2048, 0, 0),
		(drawing, 224, 0, 2048, 0, 0),
		(drawing, 225, 0, 2048, 0, 0),
		(drawing, 226, 0, 2048, 0, 0),
		(drawing, 227, 0, 2048, 0, 0),
		(drawing, 228, 0, 2048, 0, 0),
		(drawing, 229, 0, 2048, 0, 0),
		(drawing, 230, 0, 2048, 0, 0),
		(drawing, 231, 0, 2048, 0, 0),
		(drawing, 232, 0, 2048, 0, 0),
		(drawing, 233, 0, 2048, 0, 0),
		(drawing, 234, 0, 2048, 0, 0),
		(drawing, 235, 0, 2048, 0, 0),
		(drawing, 236, 0, 2048, 0, 0),
		(drawing, 237, 0, 2048, 0, 0),
		(drawing, 238, 0, 2048, 0, 0),
		(drawing, 239, 0, 2048, 0, 0),
		(drawing, 240, 0, 2048, 0, 0),
		(drawing, 241, 0, 2048, 0, 0),
		(drawing, 242, 0, 2048, 0, 0),
		(drawing, 243, 0, 2048, 0, 0),
		(drawing, 244, 0, 2048, 0, 0),
		(drawing, 245, 0, 2048, 0, 0),
		(drawing, 246, 0, 2048, 0, 0),
		(drawing, 247, 0, 2048, 0, 0),
		(drawing, 248, 0, 2048, 0, 0),
		(drawing, 249, 0, 2048, 0, 0),
		(drawing, 250, 0, 2048, 0, 0),
		(drawing, 251, 0, 2048, 0, 0),
		(drawing, 252, 0, 2048, 0, 0),
		(drawing, 253, 0, 2048, 0, 0),
		(drawing, 254, 0, 2048, 0, 0),
		(drawing, 255, 0, 2048, 0, 0),
		(drawing, 256, 0, 2048, 0, 0),
		(drawing, 257, 0, 2048, 0, 0),
		(drawing, 258, 0, 2048, 0, 0),
		(drawing, 259, 0, 2048, 0, 0),
		(drawing, 260, 0, 2048, 0, 0),
		(drawing, 261, 0, 2048, 0, 0),
		(drawing, 262, 0, 2048, 0, 0),
		(drawing, 263, 0, 2048, 0, 0),
		(drawing, 264, 0, 2048, 0, 0),
		(drawing, 265, 0, 2048, 0, 0),
		(drawing, 266, 0, 2048, 0, 0),
		(drawing, 267, 0, 2048, 0, 0),
		(drawing, 268, 0, 2048, 0, 0),
		(drawing, 269, 0, 2048, 0, 0),
		(drawing, 270, 0, 2048, 0, 0),
		(drawing, 271, 0, 2048, 0, 0),
		(drawing, 272, 0, 2048, 0, 0),
		(drawing, 273, 0, 2048, 0, 0),
		(drawing, 274, 0, 2048, 0, 0),
		(drawing, 275, 0, 2048, 0, 0),
		(drawing, 276, 0, 2048, 0, 0),
		(drawing, 277, 0, 2048, 0, 0),
		(drawing, 278, 0, 2048, 0, 0),
		(drawing, 279, 0, 2048, 0, 0),
		(drawing, 280, 0, 2048, 0, 0),
		(drawing, 281, 0, 2048, 0, 0),
		(drawing, 282, 0, 2048, 0, 0),
		(drawing, 283, 0, 2048, 0, 0),
		(drawing, 284, 0, 2048, 0, 0),
		(drawing, 285, 0, 2048, 0, 0),
		(drawing, 286, 0, 2048, 0, 0),
		(drawing, 287, 0, 2048, 0, 0),
		(drawing, 288, 0, 2048, 0, 0),
		(drawing, 289, 0, 2048, 0, 0),
		(drawing, 290, 0, 2048, 0, 0),
		(drawing, 291, 0, 2048, 0, 0),
		(drawing, 292, 0, 2048, 0, 0),
		(drawing, 293, 0, 2048, 0, 0),
		(drawing, 294, 0, 2048, 0, 0),
		(drawing, 295, 0, 2048, 0, 0),
		(drawing, 296, 0, 2048, 0, 0),
		(drawing, 297, 0, 2048, 0, 0),
		(drawing, 298, 0, 2048, 0, 0),
		(drawing, 299, 0, 2048, 0, 0),
		(drawing, 300, 0, 2048, 0, 0),
		(drawing, 301, 0, 2048, 0, 0),
		(drawing, 302, 0, 2048, 0, 0),
		(drawing, 303, 0, 2048, 0, 0),
		(drawing, 304, 0, 2048, 0, 0),
		(drawing, 305, 0, 2048, 0, 0),
		(drawing, 306, 0, 2048, 0, 0),
		(drawing, 307, 0, 2048, 0, 0),
		(drawing, 308, 0, 2048, 0, 0),
		(drawing, 309, 0, 2048, 0, 0),
		(drawing, 310, 0, 2048, 0, 0),
		(drawing, 311, 0, 2048, 0, 0),
		(drawing, 312, 0, 2048, 0, 0),
		(drawing, 313, 0, 2048, 0, 0),
		(drawing, 314, 0, 2048, 0, 0),
		(drawing, 315, 0, 2048, 0, 0),
		(drawing, 316, 0, 2048, 0, 0),
		(drawing, 317, 0, 2048, 0, 0),
		(drawing, 318, 0, 2048, 0, 0),
		(drawing, 319, 0, 2048, 0, 0),
		(drawing, 320, 0, 2048, 0, 0),
		(drawing, 321, 0, 2048, 0, 0),
		(drawing, 322, 0, 2048, 0, 0),
		(drawing, 323, 0, 2048, 0, 0),
		(drawing, 324, 0, 2048, 0, 0),
		(drawing, 325, 0, 2048, 0, 0),
		(drawing, 326, 0, 2048, 0, 0),
		(drawing, 327, 0, 2048, 0, 0),
		(drawing, 328, 0, 2048, 0, 0),
		(drawing, 329, 0, 2048, 0, 0),
		(drawing, 330, 0, 2048, 0, 0),
		(drawing, 331, 0, 2048, 0, 0),
		(drawing, 332, 0, 2048, 0, 0),
		(drawing, 333, 0, 2048, 0, 0),
		(drawing, 334, 0, 2048, 0, 0),
		(drawing, 335, 0, 2048, 0, 0),
		(drawing, 336, 0, 2048, 0, 0),
		(drawing, 337, 0, 2048, 0, 0),
		(drawing, 338, 0, 2048, 0, 0),
		(drawing, 339, 0, 2048, 0, 0),
		(drawing, 340, 0, 2048, 0, 0),
		(drawing, 341, 0, 2048, 0, 0),
		(drawing, 342, 0, 2048, 0, 0),
		(drawing, 343, 0, 2048, 0, 0),
		(drawing, 344, 0, 2048, 0, 0),
		(drawing, 345, 0, 2048, 0, 0),
		(drawing, 346, 0, 2048, 0, 0),
		(drawing, 347, 0, 2048, 0, 0),
		(drawing, 348, 0, 2048, 0, 0),
		(drawing, 349, 0, 2048, 0, 0),
		(drawing, 350, 0, 2048, 0, 0),
		(drawing, 351, 0, 2048, 0, 0),
		(drawing, 352, 0, 2048, 0, 0),
		(drawing, 353, 0, 2048, 0, 0),
		(drawing, 354, 0, 2048, 0, 0),
		(drawing, 355, 0, 2048, 0, 0),
		(drawing, 356, 0, 2048, 0, 0),
		(drawing, 357, 0, 2048, 0, 0),
		(drawing, 358, 0, 2048, 0, 0),
		(drawing, 359, 0, 2048, 0, 0),
		(drawing, 360, 0, 2048, 0, 0),
		(drawing, 361, 0, 2048, 0, 0),
		(drawing, 362, 0, 2048, 0, 0),
		(drawing, 363, 0, 2048, 0, 0),
		(drawing, 364, 0, 2048, 0, 0),
		(drawing, 365, 0, 2048, 0, 0),
		(drawing, 366, 0, 2048, 0, 0),
		(drawing, 367, 0, 2048, 0, 0),
		(drawing, 368, 0, 2048, 0, 0),
		(drawing, 369, 0, 2048, 0, 0),
		(drawing, 370, 0, 2048, 0, 0),
		(drawing, 371, 0, 2048, 0, 0),
		(drawing, 372, 0, 2048, 0, 0),
		(drawing, 373, 0, 2048, 0, 0),
		(drawing, 374, 0, 2048, 0, 0),
		(drawing, 375, 0, 2048, 0, 0),
		(drawing, 376, 0, 2048, 0, 0),
		(drawing, 377, 0, 2048, 0, 0),
		(drawing, 378, 0, 2048, 0, 0),
		(drawing, 379, 0, 2048, 0, 0),
		(drawing, 380, 0, 2048, 0, 0),
		(drawing, 381, 0, 2048, 0, 0),
		(drawing, 382, 0, 2048, 0, 0),
		(drawing, 383, 0, 2048, 0, 0),
		(drawing, 384, 0, 2048, 0, 0),
		(drawing, 385, 0, 2048, 0, 0),
		(drawing, 386, 0, 2048, 0, 0),
		(drawing, 387, 0, 2048, 0, 0),
		(drawing, 388, 0, 2048, 0, 0),
		(drawing, 389, 0, 2048, 0, 0),
		(drawing, 390, 0, 2048, 0, 0),
		(drawing, 391, 0, 2048, 0, 0),
		(drawing, 392, 0, 2048, 0, 0),
		(drawing, 393, 0, 2048, 0, 0),
		(drawing, 394, 0, 2048, 0, 0),
		(drawing, 395, 0, 2048, 0, 0),
		(drawing, 396, 0, 2048, 0, 0),
		(drawing, 397, 0, 2048, 0, 0),
		(drawing, 398, 0, 2048, 0, 0),
		(drawing, 399, 0, 2048, 0, 0),
		(drawing, 400, 0, 2048, 0, 0),
		(drawing, 401, 0, 2048, 0, 0),
		(drawing, 402, 0, 2048, 0, 0),
		(drawing, 403, 0, 2048, 0, 0),
		(drawing, 404, 0, 2048, 0, 0),
		(drawing, 405, 0, 2048, 0, 0),
		(drawing, 406, 0, 2048, 0, 0),
		(drawing, 407, 0, 2048, 0, 0),
		(drawing, 408, 0, 2048, 0, 0),
		(drawing, 409, 0, 2048, 0, 0),
		(drawing, 410, 0, 2048, 0, 0),
		(drawing, 411, 0, 2048, 0, 0),
		(drawing, 412, 0, 2048, 0, 0),
		(drawing, 413, 0, 2048, 0, 0),
		(drawing, 414, 0, 2048, 0, 0),
		(drawing, 415, 0, 2048, 0, 0),
		(drawing, 416, 0, 2048, 0, 0),
		(drawing, 417, 0, 2048, 0, 0),
		(drawing, 418, 0, 2048, 0, 0),
		(drawing, 419, 0, 2048, 0, 0),
		(drawing, 420, 0, 2048, 0, 0),
		(drawing, 421, 0, 2048, 0, 0),
		(drawing, 422, 0, 2048, 0, 0),
		(drawing, 423, 0, 2048, 0, 0),
		(drawing, 424, 0, 2048, 0, 0),
		(drawing, 425, 0, 2048, 0, 0),
		(drawing, 426, 0, 2048, 0, 0),
		(drawing, 427, 0, 2048, 0, 0),
		(drawing, 428, 0, 2048, 0, 0),
		(drawing, 429, 0, 2048, 0, 0),
		(drawing, 430, 0, 2048, 0, 0),
		(drawing, 431, 0, 2048, 0, 0),
		(drawing, 432, 0, 2048, 0, 0),
		(drawing, 433, 0, 2048, 0, 0),
		(drawing, 434, 0, 2048, 0, 0),
		(drawing, 435, 0, 2048, 0, 0),
		(drawing, 436, 0, 2048, 0, 0),
		(drawing, 437, 0, 2048, 0, 0),
		(drawing, 438, 0, 2048, 0, 0),
		(drawing, 439, 0, 2048, 0, 0),
		(drawing, 440, 0, 2048, 0, 0),
		(drawing, 441, 0, 2048, 0, 0),
		(drawing, 442, 0, 2048, 0, 0),
		(drawing, 443, 0, 2048, 0, 0),
		(drawing, 444, 0, 2048, 0, 0),
		(drawing, 445, 0, 2048, 0, 0),
		(drawing, 446, 0, 2048, 0, 0),
		(drawing, 447, 0, 2048, 0, 0),
		(drawing, 448, 0, 2048, 0, 0),
		(drawing, 449, 0, 2048, 0, 0),
		(drawing, 450, 0, 2048, 0, 0),
		(drawing, 451, 0, 2048, 0, 0),
		(drawing, 452, 0, 2048, 0, 0),
		(drawing, 453, 0, 2048, 0, 0),
		(drawing, 454, 0, 2048, 0, 0),
		(drawing, 455, 0, 2048, 0, 0),
		(drawing, 456, 0, 2048, 0, 0),
		(drawing, 457, 0, 2048, 0, 0),
		(drawing, 458, 0, 2048, 0, 0),
		(drawing, 459, 0, 2048, 0, 0),
		(drawing, 460, 0, 2048, 0, 0),
		(drawing, 461, 0, 2048, 0, 0),
		(drawing, 462, 0, 2048, 0, 0),
		(drawing, 463, 0, 2048, 0, 0),
		(drawing, 464, 0, 2048, 0, 0),
		(drawing, 465, 0, 2048, 0, 0),
		(drawing, 466, 0, 2048, 0, 0),
		(drawing, 467, 0, 2048, 0, 0),
		(drawing, 468, 0, 2048, 0, 0),
		(drawing, 469, 0, 2048, 0, 0),
		(drawing, 470, 0, 2048, 0, 0),
		(drawing, 471, 0, 2048, 0, 0),
		(drawing, 472, 0, 2048, 0, 0),
		(drawing, 473, 0, 2048, 0, 0),
		(drawing, 474, 0, 2048, 0, 0),
		(drawing, 475, 0, 2048, 0, 0),
		(drawing, 476, 0, 2048, 0, 0),
		(drawing, 477, 0, 2048, 0, 0),
		(drawing, 478, 0, 2048, 0, 0),
		(drawing, 479, 0, 2048, 0, 0),
		(drawing, 480, 0, 2048, 0, 0),
		(drawing, 481, 0, 2048, 0, 0),
		(drawing, 482, 0, 2048, 0, 0),
		(drawing, 483, 0, 2048, 0, 0),
		(drawing, 484, 0, 2048, 0, 0),
		(drawing, 485, 0, 2048, 0, 0),
		(drawing, 486, 0, 2048, 0, 0),
		(drawing, 487, 0, 2048, 0, 0),
		(drawing, 488, 0, 2048, 0, 0),
		(drawing, 489, 0, 2048, 0, 0),
		(drawing, 490, 0, 2048, 0, 0),
		(drawing, 491, 0, 2048, 0, 0),
		(drawing, 492, 0, 2048, 0, 0),
		(drawing, 493, 0, 2048, 0, 0),
		(drawing, 494, 0, 2048, 0, 0),
		(drawing, 495, 0, 2048, 0, 0),
		(drawing, 496, 0, 2048, 0, 0),
		(drawing, 497, 0, 2048, 0, 0),
		(drawing, 498, 0, 2048, 0, 0),
		(drawing, 499, 0, 2048, 0, 0),
		(drawing, 500, 0, 2048, 0, 0),
		(drawing, 501, 0, 2048, 0, 0),
		(drawing, 502, 0, 2048, 0, 0),
		(drawing, 503, 0, 2048, 0, 0),
		(drawing, 504, 0, 2048, 0, 0),
		(drawing, 505, 0, 2048, 0, 0),
		(drawing, 506, 0, 2048, 0, 0),
		(drawing, 507, 0, 2048, 0, 0),
		(drawing, 508, 0, 2048, 0, 0),
		(drawing, 509, 0, 2048, 0, 0),
		(drawing, 510, 0, 2048, 0, 0),
		(drawing, 511, 0, 2048, 0, 0),
		(drawing, 512, 0, 2048, 0, 0),
		(drawing, 513, 0, 2048, 0, 0),
		(drawing, 514, 0, 2048, 0, 0),
		(drawing, 515, 0, 2048, 0, 0),
		(drawing, 516, 0, 2048, 0, 0),
		(drawing, 517, 0, 2048, 0, 0),
		(drawing, 518, 0, 2048, 0, 0),
		(drawing, 519, 0, 2048, 0, 0),
		(drawing, 520, 0, 2048, 0, 0),
		(drawing, 521, 0, 2048, 0, 0),
		(drawing, 522, 0, 2048, 0, 0),
		(drawing, 523, 0, 2048, 0, 0),
		(drawing, 524, 0, 2048, 0, 0),
		(drawing, 525, 0, 2048, 0, 0),
		(drawing, 526, 0, 2048, 0, 0),
		(drawing, 527, 0, 2048, 0, 0),
		(drawing, 528, 0, 2048, 0, 0),
		(drawing, 529, 0, 2048, 0, 0),
		(drawing, 530, 0, 2048, 0, 0),
		(drawing, 531, 0, 2048, 0, 0),
		(drawing, 532, 0, 2048, 0, 0),
		(drawing, 533, 0, 2048, 0, 0),
		(drawing, 534, 0, 2048, 0, 0),
		(drawing, 535, 0, 2048, 0, 0),
		(drawing, 536, 0, 2048, 0, 0),
		(drawing, 537, 0, 2048, 0, 0),
		(drawing, 538, 0, 2048, 0, 0),
		(drawing, 539, 0, 2048, 0, 0),
		(drawing, 540, 0, 2048, 0, 0),
		(drawing, 541, 0, 2048, 0, 0),
		(drawing, 542, 0, 2048, 0, 0),
		(drawing, 543, 0, 2048, 0, 0),
		(drawing, 544, 0, 2048, 0, 0),
		(drawing, 545, 0, 2048, 0, 0),
		(drawing, 546, 0, 2048, 0, 0),
		(drawing, 547, 0, 2048, 0, 0),
		(drawing, 548, 0, 2048, 0, 0),
		(drawing, 549, 0, 2048, 0, 0),
		(drawing, 550, 0, 2048, 0, 0),
		(drawing, 551, 0, 2048, 0, 0),
		(drawing, 552, 0, 2048, 0, 0),
		(drawing, 553, 0, 2048, 0, 0),
		(drawing, 554, 0, 2048, 0, 0),
		(drawing, 555, 0, 2048, 0, 0),
		(drawing, 556, 0, 2048, 0, 0),
		(drawing, 557, 0, 2048, 0, 0),
		(drawing, 558, 0, 2048, 0, 0),
		(drawing, 559, 0, 2048, 0, 0),
		(drawing, 560, 0, 2048, 0, 0),
		(drawing, 561, 0, 2048, 0, 0),
		(drawing, 562, 0, 2048, 0, 0),
		(drawing, 563, 0, 2048, 0, 0),
		(drawing, 564, 0, 2048, 0, 0),
		(drawing, 565, 0, 2048, 0, 0),
		(drawing, 566, 0, 2048, 0, 0),
		(drawing, 567, 0, 2048, 0, 0),
		(drawing, 568, 0, 2048, 0, 0),
		(drawing, 569, 0, 2048, 0, 0),
		(drawing, 570, 0, 2048, 0, 0),
		(drawing, 571, 0, 2048, 0, 0),
		(drawing, 572, 0, 2048, 0, 0),
		(drawing, 573, 0, 2048, 0, 0),
		(drawing, 574, 0, 2048, 0, 0),
		(drawing, 575, 0, 2048, 0, 0),
		(drawing, 576, 0, 2048, 0, 0),
		(drawing, 577, 0, 2048, 0, 0),
		(drawing, 578, 0, 2048, 0, 0),
		(drawing, 579, 0, 2048, 0, 0),
		(drawing, 580, 0, 2048, 0, 0),
		(drawing, 581, 0, 2048, 0, 0),
		(drawing, 582, 0, 2048, 0, 0),
		(drawing, 583, 0, 2048, 0, 0),
		(drawing, 584, 0, 2048, 0, 0),
		(drawing, 585, 0, 2048, 0, 0),
		(drawing, 586, 0, 2048, 0, 0),
		(drawing, 587, 0, 2048, 0, 0),
		(drawing, 588, 0, 2048, 0, 0),
		(drawing, 589, 0, 2048, 0, 0),
		(drawing, 590, 0, 2048, 0, 0),
		(drawing, 591, 0, 2048, 0, 0),
		(drawing, 592, 0, 2048, 0, 0),
		(drawing, 593, 0, 2048, 0, 0),
		(drawing, 594, 0, 2048, 0, 0),
		(drawing, 595, 0, 2048, 0, 0),
		(drawing, 596, 0, 2048, 0, 0),
		(drawing, 597, 0, 2048, 0, 0),
		(drawing, 598, 0, 2048, 0, 0),
		(drawing, 599, 0, 2048, 0, 0),
		(drawing, 600, 0, 2048, 0, 0),
		(drawing, 601, 0, 2048, 0, 0),
		(drawing, 602, 0, 2048, 0, 0),
		(drawing, 603, 0, 2048, 0, 0),
		(drawing, 604, 0, 2048, 0, 0),
		(drawing, 605, 0, 2048, 0, 0),
		(drawing, 606, 0, 2048, 0, 0),
		(drawing, 607, 0, 2048, 0, 0),
		(drawing, 608, 0, 2048, 0, 0),
		(drawing, 609, 0, 2048, 0, 0),
		(drawing, 610, 0, 2048, 0, 0),
		(drawing, 611, 0, 2048, 0, 0),
		(drawing, 612, 0, 2048, 0, 0),
		(drawing, 613, 0, 2048, 0, 0),
		(drawing, 614, 0, 2048, 0, 0),
		(drawing, 615, 0, 2048, 0, 0),
		(drawing, 616, 0, 2048, 0, 0),
		(drawing, 617, 0, 2048, 0, 0),
		(drawing, 618, 0, 2048, 0, 0),
		(drawing, 619, 0, 2048, 0, 0),
		(drawing, 620, 0, 2048, 0, 0),
		(drawing, 621, 0, 2048, 0, 0),
		(drawing, 622, 0, 2048, 0, 0),
		(drawing, 623, 0, 2048, 0, 0),
		(drawing, 624, 0, 2048, 0, 0),
		(drawing, 625, 0, 2048, 0, 0),
		(drawing, 626, 0, 2048, 0, 0),
		(drawing, 627, 0, 2048, 0, 0),
		(drawing, 628, 0, 2048, 0, 0),
		(drawing, 629, 0, 2048, 0, 0),
		(drawing, 630, 0, 2048, 0, 0),
		(drawing, 631, 0, 2048, 0, 0),
		(drawing, 632, 0, 2048, 0, 0),
		(drawing, 633, 0, 2048, 0, 0),
		(drawing, 634, 0, 2048, 0, 0),
		(drawing, 635, 0, 2048, 0, 0),
		(drawing, 636, 0, 2048, 0, 0),
		(drawing, 637, 0, 2048, 0, 0),
		(drawing, 638, 0, 2048, 0, 0),
		(drawing, 639, 0, 2048, 0, 0),
		(drawing, 640, 0, 2048, 0, 0),
		(drawing, 641, 0, 2048, 0, 0),
		(drawing, 642, 0, 2048, 0, 0),
		(drawing, 643, 0, 2048, 0, 0),
		(drawing, 644, 0, 2048, 0, 0),
		(drawing, 645, 0, 2048, 0, 0),
		(drawing, 646, 0, 2048, 0, 0),
		(drawing, 647, 0, 2048, 0, 0),
		(drawing, 648, 0, 2048, 0, 0),
		(drawing, 649, 0, 2048, 0, 0),
		(drawing, 650, 0, 2048, 0, 0),
		(drawing, 651, 0, 2048, 0, 0),
		(drawing, 652, 0, 2048, 0, 0),
		(drawing, 653, 0, 2048, 0, 0),
		(drawing, 654, 0, 2048, 0, 0),
		(drawing, 655, 0, 2048, 0, 0),
		(drawing, 656, 0, 2048, 0, 0),
		(drawing, 657, 0, 2048, 0, 0),
		(drawing, 658, 0, 2048, 0, 0),
		(drawing, 659, 0, 2048, 0, 0),
		(drawing, 660, 0, 2048, 0, 0),
		(drawing, 661, 0, 2048, 0, 0),
		(drawing, 662, 0, 2048, 0, 0),
		(drawing, 663, 0, 2048, 0, 0),
		(drawing, 664, 0, 2048, 0, 0),
		(drawing, 665, 0, 2048, 0, 0),
		(drawing, 666, 0, 2048, 0, 0),
		(drawing, 667, 0, 2048, 0, 0),
		(drawing, 668, 0, 2048, 0, 0),
		(drawing, 669, 0, 2048, 0, 0),
		(drawing, 670, 0, 2048, 0, 0),
		(drawing, 671, 0, 2048, 0, 0),
		(drawing, 672, 0, 2048, 0, 0),
		(drawing, 673, 0, 2048, 0, 0),
		(drawing, 674, 0, 2048, 0, 0),
		(drawing, 675, 0, 2048, 0, 0),
		(drawing, 676, 0, 2048, 0, 0),
		(drawing, 677, 0, 2048, 0, 0),
		(drawing, 678, 0, 2048, 0, 0),
		(drawing, 679, 0, 2048, 0, 0),
		(drawing, 680, 0, 2048, 0, 0),
		(drawing, 681, 0, 2048, 0, 0),
		(drawing, 682, 0, 2048, 0, 0),
		(drawing, 683, 0, 2048, 0, 0),
		(drawing, 684, 0, 2048, 0, 0),
		(drawing, 685, 0, 2048, 0, 0),
		(drawing, 686, 0, 2048, 0, 0),
		(drawing, 687, 0, 2048, 0, 0),
		(drawing, 688, 0, 2048, 0, 0),
		(drawing, 689, 0, 2048, 0, 0),
		(drawing, 690, 0, 2048, 0, 0),
		(drawing, 691, 0, 2048, 0, 0),
		(drawing, 692, 0, 2048, 0, 0),
		(drawing, 693, 0, 2048, 0, 0),
		(drawing, 694, 0, 2048, 0, 0),
		(drawing, 695, 0, 2048, 0, 0),
		(drawing, 696, 0, 2048, 0, 0),
		(drawing, 697, 0, 2048, 0, 0),
		(drawing, 698, 0, 2048, 0, 0),
		(drawing, 699, 0, 2048, 0, 0),
		(drawing, 700, 0, 2048, 0, 0),
		(drawing, 701, 0, 2048, 0, 0),
		(drawing, 702, 0, 2048, 0, 0),
		(drawing, 703, 0, 2048, 0, 0),
		(drawing, 704, 0, 2048, 0, 0),
		(drawing, 705, 0, 2048, 0, 0),
		(drawing, 706, 0, 2048, 0, 0),
		(drawing, 707, 0, 2048, 0, 0),
		(drawing, 708, 0, 2048, 0, 0),
		(drawing, 709, 0, 2048, 0, 0),
		(drawing, 710, 0, 2048, 0, 0),
		(drawing, 711, 0, 2048, 0, 0),
		(drawing, 712, 0, 2048, 0, 0),
		(drawing, 713, 0, 2048, 0, 0),
		(drawing, 714, 0, 2048, 0, 0),
		(drawing, 715, 0, 2048, 0, 0),
		(drawing, 716, 0, 2048, 0, 0),
		(drawing, 717, 0, 2048, 0, 0),
		(drawing, 718, 0, 2048, 0, 0),
		(drawing, 719, 0, 2048, 0, 0),
		(drawing, 720, 0, 2048, 0, 0),
		(drawing, 721, 0, 2048, 0, 0),
		(drawing, 722, 0, 2048, 0, 0),
		(drawing, 723, 0, 2048, 0, 0),
		(drawing, 724, 0, 2048, 0, 0),
		(drawing, 725, 0, 2048, 0, 0),
		(drawing, 726, 0, 2048, 0, 0),
		(drawing, 727, 0, 2048, 0, 0),
		(drawing, 728, 0, 2048, 0, 0),
		(drawing, 729, 0, 2048, 0, 0),
		(drawing, 730, 0, 2048, 0, 0),
		(drawing, 731, 0, 2048, 0, 0),
		(drawing, 732, 0, 2048, 0, 0),
		(drawing, 733, 0, 2048, 0, 0),
		(drawing, 734, 0, 2048, 0, 0),
		(drawing, 735, 0, 2048, 0, 0),
		(drawing, 736, 0, 2048, 0, 0),
		(drawing, 737, 0, 2048, 0, 0),
		(drawing, 738, 0, 2048, 0, 0),
		(drawing, 739, 0, 2048, 0, 0),
		(drawing, 740, 0, 2048, 0, 0),
		(drawing, 741, 0, 2048, 0, 0),
		(drawing, 742, 0, 2048, 0, 0),
		(drawing, 743, 0, 2048, 0, 0),
		(drawing, 744, 0, 2048, 0, 0),
		(drawing, 745, 0, 2048, 0, 0),
		(drawing, 746, 0, 2048, 0, 0),
		(drawing, 747, 0, 2048, 0, 0),
		(drawing, 748, 0, 2048, 0, 0),
		(drawing, 749, 0, 2048, 0, 0),
		(drawing, 750, 0, 2048, 0, 0),
		(drawing, 751, 0, 2048, 0, 0),
		(drawing, 752, 0, 2048, 0, 0),
		(drawing, 753, 0, 2048, 0, 0),
		(drawing, 754, 0, 2048, 0, 0),
		(drawing, 755, 0, 2048, 0, 0),
		(drawing, 756, 0, 2048, 0, 0),
		(drawing, 757, 0, 2048, 0, 0),
		(drawing, 758, 0, 2048, 0, 0),
		(drawing, 759, 0, 2048, 0, 0),
		(drawing, 760, 0, 2048, 0, 0),
		(drawing, 761, 0, 2048, 0, 0),
		(drawing, 762, 0, 2048, 0, 0),
		(drawing, 763, 0, 2048, 0, 0),
		(drawing, 764, 0, 2048, 0, 0),
		(drawing, 765, 0, 2048, 0, 0),
		(drawing, 766, 0, 2048, 0, 0),
		(drawing, 767, 0, 2048, 0, 0),
		(drawing, 768, 0, 2048, 0, 0),
		(drawing, 769, 0, 2048, 0, 0),
		(drawing, 770, 0, 2048, 0, 0),
		(drawing, 771, 0, 2048, 0, 0),
		(drawing, 772, 0, 2048, 0, 0),
		(drawing, 773, 0, 2048, 0, 0),
		(drawing, 774, 0, 2048, 0, 0),
		(drawing, 775, 0, 2048, 0, 0),
		(drawing, 776, 0, 2048, 0, 0),
		(drawing, 777, 0, 2048, 0, 0),
		(drawing, 778, 0, 2048, 0, 0),
		(drawing, 779, 0, 2048, 0, 0),
		(drawing, 780, 0, 2048, 0, 0),
		(drawing, 781, 0, 2048, 0, 0),
		(drawing, 782, 0, 2048, 0, 0),
		(drawing, 783, 0, 2048, 0, 0),
		(drawing, 784, 0, 2048, 0, 0),
		(drawing, 785, 0, 2048, 0, 0),
		(drawing, 786, 0, 2048, 0, 0),
		(drawing, 787, 0, 2048, 0, 0),
		(drawing, 788, 0, 2048, 0, 0),
		(drawing, 789, 0, 2048, 0, 0),
		(drawing, 790, 0, 2048, 0, 0),
		(drawing, 791, 0, 2048, 0, 0),
		(drawing, 792, 0, 2048, 0, 0),
		(drawing, 793, 0, 2048, 0, 0),
		(drawing, 794, 0, 2048, 0, 0),
		(drawing, 795, 0, 2048, 0, 0),
		(drawing, 796, 0, 2048, 0, 0),
		(drawing, 797, 0, 2048, 0, 0),
		(drawing, 798, 0, 2048, 0, 0),
		(drawing, 799, 0, 2048, 0, 0),
		(drawing, 800, 0, 2048, 0, 0),
		(drawing, 801, 0, 2048, 0, 0),
		(drawing, 802, 0, 2048, 0, 0),
		(drawing, 803, 0, 2048, 0, 0),
		(drawing, 804, 0, 2048, 0, 0),
		(drawing, 805, 0, 2048, 0, 0),
		(drawing, 806, 0, 2048, 0, 0),
		(drawing, 807, 0, 2048, 0, 0),
		(drawing, 808, 0, 2048, 0, 0),
		(drawing, 809, 0, 2048, 0, 0),
		(drawing, 810, 0, 2048, 0, 0),
		(drawing, 811, 0, 2048, 0, 0),
		(drawing, 812, 0, 2048, 0, 0),
		(drawing, 813, 0, 2048, 0, 0),
		(drawing, 814, 0, 2048, 0, 0),
		(drawing, 815, 0, 2048, 0, 0),
		(drawing, 816, 0, 2048, 0, 0),
		(drawing, 817, 0, 2048, 0, 0),
		(drawing, 818, 0, 2048, 0, 0),
		(drawing, 819, 0, 2048, 0, 0),
		(drawing, 820, 0, 2048, 0, 0),
		(drawing, 821, 0, 2048, 0, 0),
		(drawing, 822, 0, 2048, 0, 0),
		(drawing, 823, 0, 2048, 0, 0),
		(drawing, 824, 0, 2048, 0, 0),
		(drawing, 825, 0, 2048, 0, 0),
		(drawing, 826, 0, 2048, 0, 0),
		(drawing, 827, 0, 2048, 0, 0),
		(drawing, 828, 0, 2048, 0, 0),
		(drawing, 829, 0, 2048, 0, 0),
		(drawing, 830, 0, 2048, 0, 0),
		(drawing, 831, 0, 2048, 0, 0),
		(drawing, 832, 0, 2048, 0, 0),
		(drawing, 833, 0, 2048, 0, 0),
		(drawing, 834, 0, 2048, 0, 0),
		(drawing, 835, 0, 2048, 0, 0),
		(drawing, 836, 0, 2048, 0, 0),
		(drawing, 837, 0, 2048, 0, 0),
		(drawing, 838, 0, 2048, 0, 0),
		(drawing, 839, 0, 2048, 0, 0),
		(drawing, 840, 0, 2048, 0, 0),
		(drawing, 841, 0, 2048, 0, 0),
		(drawing, 842, 0, 2048, 0, 0),
		(drawing, 843, 0, 2048, 0, 0),
		(drawing, 844, 0, 2048, 0, 0),
		(drawing, 845, 0, 2048, 0, 0),
		(drawing, 846, 0, 2048, 0, 0),
		(drawing, 847, 0, 2048, 0, 0),
		(drawing, 848, 0, 2048, 0, 0),
		(drawing, 849, 0, 2048, 0, 0),
		(drawing, 850, 0, 2048, 0, 0),
		(drawing, 851, 0, 2048, 0, 0),
		(drawing, 852, 0, 2048, 0, 0),
		(drawing, 853, 0, 2048, 0, 0),
		(drawing, 854, 0, 2048, 0, 0),
		(drawing, 855, 0, 2048, 0, 0),
		(drawing, 856, 0, 2048, 0, 0),
		(drawing, 857, 0, 2048, 0, 0),
		(drawing, 858, 0, 2048, 0, 0),
		(drawing, 859, 0, 2048, 0, 0),
		(drawing, 860, 0, 2048, 0, 0),
		(drawing, 861, 0, 2048, 0, 0),
		(drawing, 862, 0, 2048, 0, 0),
		(drawing, 863, 0, 2048, 0, 0),
		(drawing, 864, 0, 2048, 0, 0),
		(drawing, 865, 0, 2048, 0, 0),
		(drawing, 866, 0, 2048, 0, 0),
		(drawing, 867, 0, 2048, 0, 0),
		(drawing, 868, 0, 2048, 0, 0),
		(drawing, 869, 0, 2048, 0, 0),
		(drawing, 870, 0, 2048, 0, 0),
		(drawing, 871, 0, 2048, 0, 0),
		(drawing, 872, 0, 2048, 0, 0),
		(drawing, 873, 0, 2048, 0, 0),
		(drawing, 874, 0, 2048, 0, 0),
		(drawing, 875, 0, 2048, 0, 0),
		(drawing, 876, 0, 2048, 0, 0),
		(drawing, 877, 0, 2048, 0, 0),
		(drawing, 878, 0, 2048, 0, 0),
		(drawing, 879, 0, 2048, 0, 0),
		(drawing, 880, 0, 2048, 0, 0),
		(drawing, 881, 0, 2048, 0, 0),
		(drawing, 882, 0, 2048, 0, 0),
		(drawing, 883, 0, 2048, 0, 0),
		(drawing, 884, 0, 2048, 0, 0),
		(drawing, 885, 0, 2048, 0, 0),
		(drawing, 886, 0, 2048, 0, 0),
		(drawing, 887, 0, 2048, 0, 0),
		(drawing, 888, 0, 2048, 0, 0),
		(drawing, 889, 0, 2048, 0, 0),
		(drawing, 890, 0, 2048, 0, 0),
		(drawing, 891, 0, 2048, 0, 0),
		(drawing, 892, 0, 2048, 0, 0),
		(drawing, 893, 0, 2048, 0, 0),
		(drawing, 894, 0, 2048, 0, 0),
		(drawing, 895, 0, 2048, 0, 0),
		(drawing, 896, 0, 2048, 0, 0),
		(drawing, 897, 0, 2048, 0, 0),
		(drawing, 898, 0, 2048, 0, 0),
		(drawing, 899, 0, 2048, 0, 0),
		(drawing, 900, 0, 2048, 0, 0),
		(drawing, 901, 0, 2048, 0, 0),
		(drawing, 902, 0, 2048, 0, 0),
		(drawing, 903, 0, 2048, 0, 0),
		(drawing, 904, 0, 2048, 0, 0),
		(drawing, 905, 0, 2048, 0, 0),
		(drawing, 906, 0, 2048, 0, 0),
		(drawing, 907, 0, 2048, 0, 0),
		(drawing, 908, 0, 2048, 0, 0),
		(drawing, 909, 0, 2048, 0, 0),
		(drawing, 910, 0, 2048, 0, 0),
		(drawing, 911, 0, 2048, 0, 0),
		(drawing, 912, 0, 2048, 0, 0),
		(drawing, 913, 0, 2048, 0, 0),
		(drawing, 914, 0, 2048, 0, 0),
		(drawing, 915, 0, 2048, 0, 0),
		(drawing, 916, 0, 2048, 0, 0),
		(drawing, 917, 0, 2048, 0, 0),
		(drawing, 918, 0, 2048, 0, 0),
		(drawing, 919, 0, 2048, 0, 0),
		(drawing, 920, 0, 2048, 0, 0),
		(drawing, 921, 0, 2048, 0, 0),
		(drawing, 922, 0, 2048, 0, 0),
		(drawing, 923, 0, 2048, 0, 0),
		(drawing, 924, 0, 2048, 0, 0),
		(drawing, 925, 0, 2048, 0, 0),
		(drawing, 926, 0, 2048, 0, 0),
		(drawing, 927, 0, 2048, 0, 0),
		(drawing, 928, 0, 2048, 0, 0),
		(drawing, 929, 0, 2048, 0, 0),
		(drawing, 930, 0, 2048, 0, 0),
		(drawing, 931, 0, 2048, 0, 0),
		(drawing, 932, 0, 2048, 0, 0),
		(drawing, 933, 0, 2048, 0, 0),
		(drawing, 934, 0, 2048, 0, 0),
		(drawing, 935, 0, 2048, 0, 0),
		(drawing, 936, 0, 2048, 0, 0),
		(drawing, 937, 0, 2048, 0, 0),
		(drawing, 938, 0, 2048, 0, 0),
		(drawing, 939, 0, 2048, 0, 0),
		(drawing, 940, 0, 2048, 0, 0),
		(drawing, 941, 0, 2048, 0, 0),
		(drawing, 942, 0, 2048, 0, 0),
		(drawing, 943, 0, 2048, 0, 0),
		(drawing, 944, 0, 2048, 0, 0),
		(drawing, 945, 0, 2048, 0, 0),
		(drawing, 946, 0, 2048, 0, 0),
		(drawing, 947, 0, 2048, 0, 0),
		(drawing, 948, 0, 2048, 0, 0),
		(drawing, 949, 0, 2048, 0, 0),
		(drawing, 950, 0, 2048, 0, 0),
		(drawing, 951, 0, 2048, 0, 0),
		(drawing, 952, 0, 2048, 0, 0),
		(drawing, 953, 0, 2048, 0, 0),
		(drawing, 954, 0, 2048, 0, 0),
		(drawing, 955, 0, 2048, 0, 0),
		(drawing, 956, 0, 2048, 0, 0),
		(drawing, 957, 0, 2048, 0, 0),
		(drawing, 958, 0, 2048, 0, 0),
		(drawing, 959, 0, 2048, 0, 0),
		(drawing, 960, 0, 2048, 0, 0),
		(drawing, 961, 0, 2048, 0, 0),
		(drawing, 962, 0, 2048, 0, 0),
		(drawing, 963, 0, 2048, 0, 0),
		(drawing, 964, 0, 2048, 0, 0),
		(drawing, 965, 0, 2048, 0, 0),
		(drawing, 966, 0, 2048, 0, 0),
		(drawing, 967, 0, 2048, 0, 0),
		(drawing, 968, 0, 2048, 0, 0),
		(drawing, 969, 0, 2048, 0, 0),
		(drawing, 970, 0, 2048, 0, 0),
		(drawing, 971, 0, 2048, 0, 0),
		(drawing, 972, 0, 2048, 0, 0),
		(drawing, 973, 0, 2048, 0, 0),
		(drawing, 974, 0, 2048, 0, 0),
		(drawing, 975, 0, 2048, 0, 0),
		(drawing, 976, 0, 2048, 0, 0),
		(drawing, 977, 0, 2048, 0, 0),
		(drawing, 978, 0, 2048, 0, 0),
		(drawing, 979, 0, 2048, 0, 0),
		(drawing, 980, 0, 2048, 0, 0),
		(drawing, 981, 0, 2048, 0, 0),
		(drawing, 982, 0, 2048, 0, 0),
		(drawing, 983, 0, 2048, 0, 0),
		(drawing, 984, 0, 2048, 0, 0),
		(drawing, 985, 0, 2048, 0, 0),
		(drawing, 986, 0, 2048, 0, 0),
		(drawing, 987, 0, 2048, 0, 0),
		(drawing, 988, 0, 2048, 0, 0),
		(drawing, 989, 0, 2048, 0, 0),
		(drawing, 990, 0, 2048, 0, 0),
		(drawing, 991, 0, 2048, 0, 0),
		(drawing, 992, 0, 2048, 0, 0),
		(drawing, 993, 0, 2048, 0, 0),
		(drawing, 994, 0, 2048, 0, 0),
		(drawing, 995, 0, 2048, 0, 0),
		(drawing, 996, 0, 2048, 0, 0),
		(drawing, 997, 0, 2048, 0, 0),
		(drawing, 998, 0, 2048, 0, 0),
		(drawing, 999, 0, 2048, 0, 0),
		(drawing, 1000, 0, 2048, 0, 0),
		(drawing, 1001, 0, 2048, 0, 0),
		(drawing, 1002, 0, 2048, 0, 0),
		(drawing, 1003, 0, 2048, 0, 0),
		(drawing, 1004, 0, 2048, 0, 0),
		(drawing, 1005, 0, 2048, 0, 0),
		(drawing, 1006, 0, 2048, 0, 0),
		(drawing, 1007, 0, 2048, 0, 0),
		(drawing, 1008, 0, 2048, 0, 0),
		(drawing, 1009, 0, 2048, 0, 0),
		(drawing, 1010, 0, 2048, 0, 0),
		(drawing, 1011, 0, 2048, 0, 0),
		(drawing, 1012, 0, 2048, 0, 0),
		(drawing, 1013, 0, 2048, 0, 0),
		(drawing, 1014, 0, 2048, 0, 0),
		(drawing, 1015, 0, 2048, 0, 0),
		(drawing, 1016, 0, 2048, 0, 0),
		(drawing, 1017, 0, 2048, 0, 0),
		(drawing, 1018, 0, 2048, 0, 0),
		(drawing, 1019, 0, 2048, 0, 0),
		(drawing, 1020, 0, 2048, 0, 0),
		(drawing, 1021, 0, 2048, 0, 0),
		(drawing, 1022, 0, 2048, 0, 0),
		(drawing, 1023, 0, 2048, 0, 0),
		(drawing, 1024, 0, 2048, 0, 0),
		(drawing, 1025, 0, 2048, 0, 0),
		(drawing, 1026, 0, 2048, 0, 0),
		(drawing, 1027, 0, 2048, 0, 0),
		(drawing, 1028, 0, 2048, 0, 0),
		(drawing, 1029, 0, 2048, 0, 0),
		(drawing, 1030, 0, 2048, 0, 0),
		(drawing, 1031, 0, 2048, 0, 0),
		(drawing, 1032, 0, 2048, 0, 0),
		(drawing, 1033, 0, 2048, 0, 0),
		(drawing, 1034, 0, 2048, 0, 0),
		(drawing, 1035, 0, 2048, 0, 0),
		(drawing, 1036, 0, 2048, 0, 0),
		(drawing, 1037, 0, 2048, 0, 0),
		(drawing, 1038, 0, 2048, 0, 0),
		(drawing, 1039, 0, 2048, 0, 0),
		(drawing, 1040, 0, 2048, 0, 0),
		(drawing, 1041, 0, 2048, 0, 0),
		(drawing, 1042, 0, 2048, 0, 0),
		(drawing, 1043, 0, 2048, 0, 0),
		(drawing, 1044, 0, 2048, 0, 0),
		(drawing, 1045, 0, 2048, 0, 0),
		(drawing, 1046, 0, 2048, 0, 0),
		(drawing, 1047, 0, 2048, 0, 0),
		(drawing, 1048, 0, 2048, 0, 0),
		(drawing, 1049, 0, 2048, 0, 0),
		(drawing, 1050, 0, 2048, 0, 0),
		(drawing, 1051, 0, 2048, 0, 0),
		(drawing, 1052, 0, 2048, 0, 0),
		(drawing, 1053, 0, 2048, 0, 0),
		(drawing, 1054, 0, 2048, 0, 0),
		(drawing, 1055, 0, 2048, 0, 0),
		(drawing, 1056, 0, 2048, 0, 0),
		(drawing, 1057, 0, 2048, 0, 0),
		(drawing, 1058, 0, 2048, 0, 0),
		(drawing, 1059, 0, 2048, 0, 0),
		(drawing, 1060, 0, 2048, 0, 0),
		(drawing, 1061, 0, 2048, 0, 0),
		(drawing, 1062, 0, 2048, 0, 0),
		(drawing, 1063, 0, 2048, 0, 0),
		(drawing, 1064, 0, 2048, 0, 0),
		(drawing, 1065, 0, 2048, 0, 0),
		(drawing, 1066, 0, 2048, 0, 0),
		(drawing, 1067, 0, 2048, 0, 0),
		(drawing, 1068, 0, 2048, 0, 0),
		(drawing, 1069, 0, 2048, 0, 0),
		(drawing, 1070, 0, 2048, 0, 0),
		(drawing, 1071, 0, 2048, 0, 0),
		(drawing, 1072, 0, 2048, 0, 0),
		(drawing, 1073, 0, 2048, 0, 0),
		(drawing, 1074, 0, 2048, 0, 0),
		(drawing, 1075, 0, 2048, 0, 0),
		(drawing, 1076, 0, 2048, 0, 0),
		(drawing, 1077, 0, 2048, 0, 0),
		(drawing, 1078, 0, 2048, 0, 0),
		(drawing, 1079, 0, 2048, 0, 0),
		(drawing, 1080, 0, 2048, 0, 0),
		(drawing, 1081, 0, 2048, 0, 0),
		(drawing, 1082, 0, 2048, 0, 0),
		(drawing, 1083, 0, 2048, 0, 0),
		(drawing, 1084, 0, 2048, 0, 0),
		(drawing, 1085, 0, 2048, 0, 0),
		(drawing, 1086, 0, 2048, 0, 0),
		(drawing, 1087, 0, 2048, 0, 0),
		(drawing, 1088, 0, 2048, 0, 0),
		(drawing, 1089, 0, 2048, 0, 0),
		(drawing, 1090, 0, 2048, 0, 0),
		(drawing, 1091, 0, 2048, 0, 0),
		(drawing, 1092, 0, 2048, 0, 0),
		(drawing, 1093, 0, 2048, 0, 0),
		(drawing, 1094, 0, 2048, 0, 0),
		(drawing, 1095, 0, 2048, 0, 0),
		(drawing, 1096, 0, 2048, 0, 0),
		(drawing, 1097, 0, 2048, 0, 0),
		(drawing, 1098, 0, 2048, 0, 0),
		(drawing, 1099, 0, 2048, 0, 0),
		(drawing, 1100, 0, 2048, 0, 0),
		(drawing, 1101, 0, 2048, 0, 0),
		(drawing, 1102, 0, 2048, 0, 0),
		(drawing, 1103, 0, 2048, 0, 0),
		(drawing, 1104, 0, 2048, 0, 0),
		(drawing, 1105, 0, 2048, 0, 0),
		(drawing, 1106, 0, 2048, 0, 0),
		(drawing, 1107, 0, 2048, 0, 0),
		(drawing, 1108, 0, 2048, 0, 0),
		(drawing, 1109, 0, 2048, 0, 0),
		(drawing, 1110, 0, 2048, 0, 0),
		(drawing, 1111, 0, 2048, 0, 0),
		(drawing, 1112, 0, 2048, 0, 0),
		(drawing, 1113, 0, 2048, 0, 0),
		(drawing, 1114, 0, 2048, 0, 0),
		(drawing, 1115, 0, 2048, 0, 0),
		(drawing, 1116, 0, 2048, 0, 0),
		(drawing, 1117, 0, 2048, 0, 0),
		(drawing, 1118, 0, 2048, 0, 0),
		(drawing, 1119, 0, 2048, 0, 0),
		(drawing, 1120, 0, 2048, 0, 0),
		(drawing, 1121, 0, 2048, 0, 0),
		(drawing, 1122, 0, 2048, 0, 0),
		(drawing, 1123, 0, 2048, 0, 0),
		(drawing, 1124, 0, 2048, 0, 0),
		(drawing, 1125, 0, 2048, 0, 0),
		(drawing, 1126, 0, 2048, 0, 0),
		(drawing, 1127, 0, 2048, 0, 0),
		(drawing, 1128, 0, 2048, 0, 0),
		(drawing, 1129, 0, 2048, 0, 0),
		(drawing, 1130, 0, 2048, 0, 0),
		(drawing, 1131, 0, 2048, 0, 0),
		(drawing, 1132, 0, 2048, 0, 0),
		(drawing, 1133, 0, 2048, 0, 0),
		(drawing, 1134, 0, 2048, 0, 0),
		(drawing, 1135, 0, 2048, 0, 0),
		(drawing, 1136, 0, 2048, 0, 0),
		(drawing, 1137, 0, 2048, 0, 0),
		(drawing, 1138, 0, 2048, 0, 0),
		(drawing, 1139, 0, 2048, 0, 0),
		(drawing, 1140, 0, 2048, 0, 0),
		(drawing, 1141, 0, 2048, 0, 0),
		(drawing, 1142, 0, 2048, 0, 0),
		(drawing, 1143, 0, 2048, 0, 0),
		(drawing, 1144, 0, 2048, 0, 0),
		(drawing, 1145, 0, 2048, 0, 0),
		(drawing, 1146, 0, 2048, 0, 0),
		(drawing, 1147, 0, 2048, 0, 0),
		(drawing, 1148, 0, 2048, 0, 0),
		(drawing, 1149, 0, 2048, 0, 0),
		(drawing, 1150, 0, 2048, 0, 0),
		(drawing, 1151, 0, 2048, 0, 0),
		(drawing, 1152, 0, 2048, 0, 0),
		(drawing, 1153, 0, 2048, 0, 0),
		(drawing, 1154, 0, 2048, 0, 0),
		(drawing, 1155, 0, 2048, 0, 0),
		(drawing, 1156, 0, 2048, 0, 0),
		(drawing, 1157, 0, 2048, 0, 0),
		(drawing, 1158, 0, 2048, 0, 0),
		(drawing, 1159, 0, 2048, 0, 0),
		(drawing, 1160, 0, 2048, 0, 0),
		(drawing, 1161, 0, 2048, 0, 0),
		(drawing, 1162, 0, 2048, 0, 0),
		(drawing, 1163, 0, 2048, 0, 0),
		(drawing, 1164, 0, 2048, 0, 0),
		(drawing, 1165, 0, 2048, 0, 0),
		(drawing, 1166, 0, 2048, 0, 0),
		(drawing, 1167, 0, 2048, 0, 0),
		(drawing, 1168, 0, 2048, 0, 0),
		(drawing, 1169, 0, 2048, 0, 0),
		(drawing, 1170, 0, 2048, 0, 0),
		(drawing, 1171, 0, 2048, 0, 0),
		(drawing, 1172, 0, 2048, 0, 0),
		(drawing, 1173, 0, 2048, 0, 0),
		(drawing, 1174, 0, 2048, 0, 0),
		(drawing, 1175, 0, 2048, 0, 0),
		(drawing, 1176, 0, 2048, 0, 0),
		(drawing, 1177, 0, 2048, 0, 0),
		(drawing, 1178, 0, 2048, 0, 0),
		(drawing, 1179, 0, 2048, 0, 0),
		(drawing, 1180, 0, 2048, 0, 0),
		(drawing, 1181, 0, 2048, 0, 0),
		(drawing, 1182, 0, 2048, 0, 0),
		(drawing, 1183, 0, 2048, 0, 0),
		(drawing, 1184, 0, 2048, 0, 0),
		(drawing, 1185, 0, 2048, 0, 0),
		(drawing, 1186, 0, 2048, 0, 0),
		(drawing, 1187, 0, 2048, 0, 0),
		(drawing, 1188, 0, 2048, 0, 0),
		(drawing, 1189, 0, 2048, 0, 0),
		(drawing, 1190, 0, 2048, 0, 0),
		(drawing, 1191, 0, 2048, 0, 0),
		(drawing, 1192, 0, 2048, 0, 0),
		(drawing, 1193, 0, 2048, 0, 0),
		(drawing, 1194, 0, 2048, 0, 0),
		(drawing, 1195, 0, 2048, 0, 0),
		(drawing, 1196, 0, 2048, 0, 0),
		(drawing, 1197, 0, 2048, 0, 0),
		(drawing, 1198, 0, 2048, 0, 0),
		(drawing, 1199, 0, 2048, 0, 0),
		(drawing, 1200, 0, 2048, 0, 0),
		(drawing, 1201, 0, 2048, 0, 0),
		(drawing, 1202, 0, 2048, 0, 0),
		(drawing, 1203, 0, 2048, 0, 0),
		(drawing, 1204, 0, 2048, 0, 0),
		(drawing, 1205, 0, 2048, 0, 0),
		(drawing, 1206, 0, 2048, 0, 0),
		(drawing, 1207, 0, 2048, 0, 0),
		(drawing, 1208, 0, 2048, 0, 0),
		(drawing, 1209, 0, 2048, 0, 0),
		(drawing, 1210, 0, 2048, 0, 0),
		(drawing, 1211, 0, 2048, 0, 0),
		(drawing, 1212, 0, 2048, 0, 0),
		(drawing, 1213, 0, 2048, 0, 0),
		(drawing, 1214, 0, 2048, 0, 0),
		(drawing, 1215, 0, 2048, 0, 0),
		(drawing, 1216, 0, 2048, 0, 0),
		(drawing, 1217, 0, 2048, 0, 0),
		(drawing, 1218, 0, 2048, 0, 0),
		(drawing, 1219, 0, 2048, 0, 0),
		(drawing, 1220, 0, 2048, 0, 0),
		(drawing, 1221, 0, 2048, 0, 0),
		(drawing, 1222, 0, 2048, 0, 0),
		(drawing, 1223, 0, 2048, 0, 0),
		(drawing, 1224, 0, 2048, 0, 0),
		(drawing, 1225, 0, 2048, 0, 0),
		(drawing, 1226, 0, 2048, 0, 0),
		(drawing, 1227, 0, 2048, 0, 0),
		(drawing, 1228, 0, 2048, 0, 0),
		(drawing, 1229, 0, 2048, 0, 0),
		(drawing, 1230, 0, 2048, 0, 0),
		(drawing, 1231, 0, 2048, 0, 0),
		(drawing, 1232, 0, 2048, 0, 0),
		(drawing, 1233, 0, 2048, 0, 0),
		(drawing, 1234, 0, 2048, 0, 0),
		(drawing, 1235, 0, 2048, 0, 0),
		(drawing, 1236, 0, 2048, 0, 0),
		(drawing, 1237, 0, 2048, 0, 0),
		(drawing, 1238, 0, 2048, 0, 0),
		(drawing, 1239, 0, 2048, 0, 0),
		(drawing, 1240, 0, 2048, 0, 0),
		(drawing, 1241, 0, 2048, 0, 0),
		(drawing, 1242, 0, 2048, 0, 0),
		(drawing, 1243, 0, 2048, 0, 0),
		(drawing, 1244, 0, 2048, 0, 0),
		(drawing, 1245, 0, 2048, 0, 0),
		(drawing, 1246, 0, 2048, 0, 0),
		(drawing, 1247, 0, 2048, 0, 0),
		(drawing, 1248, 0, 2048, 0, 0),
		(drawing, 1249, 0, 2048, 0, 0),
		(drawing, 1250, 0, 2048, 0, 0),
		(drawing, 1251, 0, 2048, 0, 0),
		(drawing, 1252, 0, 2048, 0, 0),
		(drawing, 1253, 0, 2048, 0, 0),
		(drawing, 1254, 0, 2048, 0, 0),
		(drawing, 1255, 0, 2048, 0, 0),
		(drawing, 1256, 0, 2048, 0, 0),
		(drawing, 1257, 0, 2048, 0, 0),
		(drawing, 1258, 0, 2048, 0, 0),
		(drawing, 1259, 0, 2048, 0, 0),
		(drawing, 1260, 0, 2048, 0, 0),
		(drawing, 1261, 0, 2048, 0, 0),
		(drawing, 1262, 0, 2048, 0, 0),
		(drawing, 1263, 0, 2048, 0, 0),
		(drawing, 1264, 0, 2048, 0, 0),
		(drawing, 1265, 0, 2048, 0, 0),
		(drawing, 1266, 0, 2048, 0, 0),
		(drawing, 1267, 0, 2048, 0, 0),
		(drawing, 1268, 0, 2048, 0, 0),
		(drawing, 1269, 0, 2048, 0, 0),
		(drawing, 1270, 0, 2048, 0, 0),
		(drawing, 1271, 0, 2048, 0, 0),
		(drawing, 1272, 0, 2048, 0, 0),
		(drawing, 1273, 0, 2048, 0, 0),
		(drawing, 1274, 0, 2048, 0, 0),
		(drawing, 1275, 0, 2048, 0, 0),
		(drawing, 1276, 0, 2048, 0, 0),
		(drawing, 1277, 0, 2048, 0, 0),
		(drawing, 1278, 0, 2048, 0, 0),
		(drawing, 1279, 0, 2048, 0, 0),
		(drawing, 1280, 0, 2048, 0, 0),
		(drawing, 1281, 0, 2048, 0, 0),
		(drawing, 1282, 0, 2048, 0, 0),
		(drawing, 1283, 0, 2048, 0, 0),
		(drawing, 1284, 0, 2048, 0, 0),
		(drawing, 1285, 0, 2048, 0, 0),
		(drawing, 1286, 0, 2048, 0, 0),
		(drawing, 1287, 0, 2048, 0, 0),
		(drawing, 1288, 0, 2048, 0, 0),
		(drawing, 1289, 0, 2048, 0, 0),
		(drawing, 1290, 0, 2048, 0, 0),
		(drawing, 1291, 0, 2048, 0, 0),
		(drawing, 1292, 0, 2048, 0, 0),
		(drawing, 1293, 0, 2048, 0, 0),
		(drawing, 1294, 0, 2048, 0, 0),
		(drawing, 1295, 0, 2048, 0, 0),
		(drawing, 1296, 0, 2048, 0, 0),
		(drawing, 1297, 0, 2048, 0, 0),
		(drawing, 1298, 0, 2048, 0, 0),
		(drawing, 1299, 0, 2048, 0, 0),
		(drawing, 1300, 0, 2048, 0, 0),
		(drawing, 1301, 0, 2048, 0, 0),
		(drawing, 1302, 0, 2048, 0, 0),
		(drawing, 1303, 0, 2048, 0, 0),
		(drawing, 1304, 0, 2048, 0, 0),
		(drawing, 1305, 0, 2048, 0, 0),
		(drawing, 1306, 0, 2048, 0, 0),
		(drawing, 1307, 0, 2048, 0, 0),
		(drawing, 1308, 0, 2048, 0, 0),
		(drawing, 1309, 0, 2048, 0, 0),
		(drawing, 1310, 0, 2048, 0, 0),
		(drawing, 1311, 0, 2048, 0, 0),
		(drawing, 1312, 0, 2048, 0, 0),
		(drawing, 1313, 0, 2048, 0, 0),
		(drawing, 1314, 0, 2048, 0, 0),
		(drawing, 1315, 0, 2048, 0, 0),
		(drawing, 1316, 0, 2048, 0, 0),
		(drawing, 1317, 0, 2048, 0, 0),
		(drawing, 1318, 0, 2048, 0, 0),
		(drawing, 1319, 0, 2048, 0, 0),
		(drawing, 1320, 0, 2048, 0, 0),
		(drawing, 1321, 0, 2048, 0, 0),
		(drawing, 1322, 0, 2048, 0, 0),
		(drawing, 1323, 0, 2048, 0, 0),
		(drawing, 1324, 0, 2048, 0, 0),
		(drawing, 1325, 0, 2048, 0, 0),
		(drawing, 1326, 0, 2048, 0, 0),
		(drawing, 1327, 0, 2048, 0, 0),
		(drawing, 1328, 0, 2048, 0, 0),
		(drawing, 1329, 0, 2048, 0, 0),
		(drawing, 1330, 0, 2048, 0, 0),
		(drawing, 1331, 0, 2048, 0, 0),
		(drawing, 1332, 0, 2048, 0, 0),
		(drawing, 1333, 0, 2048, 0, 0),
		(drawing, 1334, 0, 2048, 0, 0),
		(drawing, 1335, 0, 2048, 0, 0),
		(drawing, 1336, 0, 2048, 0, 0),
		(drawing, 1337, 0, 2048, 0, 0),
		(drawing, 1338, 0, 2048, 0, 0),
		(drawing, 1339, 0, 2048, 0, 0),
		(drawing, 1340, 0, 2048, 0, 0),
		(drawing, 1341, 0, 2048, 0, 0),
		(drawing, 1342, 0, 2048, 0, 0),
		(drawing, 1343, 0, 2048, 0, 0),
		(drawing, 1344, 0, 2048, 0, 0),
		(drawing, 1345, 0, 2048, 0, 0),
		(drawing, 1346, 0, 2048, 0, 0),
		(drawing, 1347, 0, 2048, 0, 0),
		(drawing, 1348, 0, 2048, 0, 0),
		(drawing, 1349, 0, 2048, 0, 0),
		(drawing, 1350, 0, 2048, 0, 0),
		(drawing, 1351, 0, 2048, 0, 0),
		(drawing, 1352, 0, 2048, 0, 0),
		(drawing, 1353, 0, 2048, 0, 0),
		(drawing, 1354, 0, 2048, 0, 0),
		(drawing, 1355, 0, 2048, 0, 0),
		(drawing, 1356, 0, 2048, 0, 0),
		(drawing, 1357, 0, 2048, 0, 0),
		(drawing, 1358, 0, 2048, 0, 0),
		(drawing, 1359, 0, 2048, 0, 0),
		(drawing, 1360, 0, 2048, 0, 0),
		(drawing, 1361, 0, 2048, 0, 0),
		(drawing, 1362, 0, 2048, 0, 0),
		(drawing, 1363, 0, 2048, 0, 0),
		(drawing, 1364, 0, 2048, 0, 0),
		(drawing, 1365, 0, 2048, 0, 0),
		(drawing, 1366, 0, 2048, 0, 0),
		(drawing, 1367, 0, 2048, 0, 0),
		(drawing, 1368, 0, 2048, 0, 0),
		(drawing, 1369, 0, 2048, 0, 0),
		(drawing, 1370, 0, 2048, 0, 0),
		(drawing, 1371, 0, 2048, 0, 0),
		(drawing, 1372, 0, 2048, 0, 0),
		(drawing, 1373, 0, 2048, 0, 0),
		(drawing, 1374, 0, 2048, 0, 0),
		(drawing, 1375, 0, 2048, 0, 0),
		(drawing, 1376, 0, 2048, 0, 0),
		(drawing, 1377, 0, 2048, 0, 0),
		(drawing, 1378, 0, 2048, 0, 0),
		(drawing, 1379, 0, 2048, 0, 0),
		(drawing, 1380, 0, 2048, 0, 0),
		(drawing, 1381, 0, 2048, 0, 0),
		(drawing, 1382, 0, 2048, 0, 0),
		(drawing, 1383, 0, 2048, 0, 0),
		(drawing, 1384, 0, 2048, 0, 0),
		(drawing, 1385, 0, 2048, 0, 0),
		(drawing, 1386, 0, 2048, 0, 0),
		(drawing, 1387, 0, 2048, 0, 0),
		(drawing, 1388, 0, 2048, 0, 0),
		(drawing, 1389, 0, 2048, 0, 0),
		(drawing, 1390, 0, 2048, 0, 0),
		(drawing, 1391, 0, 2048, 0, 0),
		(drawing, 1392, 0, 2048, 0, 0),
		(drawing, 1393, 0, 2048, 0, 0),
		(drawing, 1394, 0, 2048, 0, 0),
		(drawing, 1395, 0, 2048, 0, 0),
		(drawing, 1396, 0, 2048, 0, 0),
		(drawing, 1397, 0, 2048, 0, 0),
		(drawing, 1398, 0, 2048, 0, 0),
		(drawing, 1399, 0, 2048, 0, 0),
		(drawing, 1400, 0, 2048, 0, 0),
		(drawing, 1401, 0, 2048, 0, 0),
		(drawing, 1402, 0, 2048, 0, 0),
		(drawing, 1403, 0, 2048, 0, 0),
		(drawing, 1404, 0, 2048, 0, 0),
		(drawing, 1405, 0, 2048, 0, 0),
		(drawing, 1406, 0, 2048, 0, 0),
		(drawing, 1407, 0, 2048, 0, 0),
		(drawing, 1408, 0, 2048, 0, 0),
		(drawing, 1409, 0, 2048, 0, 0),
		(drawing, 1410, 0, 2048, 0, 0),
		(drawing, 1411, 0, 2048, 0, 0),
		(drawing, 1412, 0, 2048, 0, 0),
		(drawing, 1413, 0, 2048, 0, 0),
		(drawing, 1414, 0, 2048, 0, 0),
		(drawing, 1415, 0, 2048, 0, 0),
		(drawing, 1416, 0, 2048, 0, 0),
		(drawing, 1417, 0, 2048, 0, 0),
		(drawing, 1418, 0, 2048, 0, 0),
		(drawing, 1419, 0, 2048, 0, 0),
		(drawing, 1420, 0, 2048, 0, 0),
		(drawing, 1421, 0, 2048, 0, 0),
		(drawing, 1422, 0, 2048, 0, 0),
		(drawing, 1423, 0, 2048, 0, 0),
		(drawing, 1424, 0, 2048, 0, 0),
		(drawing, 1425, 0, 2048, 0, 0),
		(drawing, 1426, 0, 2048, 0, 0),
		(drawing, 1427, 0, 2048, 0, 0),
		(drawing, 1428, 0, 2048, 0, 0),
		(drawing, 1429, 0, 2048, 0, 0),
		(drawing, 1430, 0, 2048, 0, 0),
		(drawing, 1431, 0, 2048, 0, 0),
		(drawing, 1432, 0, 2048, 0, 0),
		(drawing, 1433, 0, 2048, 0, 0),
		(drawing, 1434, 0, 2048, 0, 0),
		(drawing, 1435, 0, 2048, 0, 0),
		(drawing, 1436, 0, 2048, 0, 0),
		(drawing, 1437, 0, 2048, 0, 0),
		(drawing, 1438, 0, 2048, 0, 0),
		(drawing, 1439, 0, 2048, 0, 0),
		(drawing, 1440, 0, 2048, 0, 0),
		(drawing, 1441, 0, 2048, 0, 0),
		(drawing, 1442, 0, 2048, 0, 0),
		(drawing, 1443, 0, 2048, 0, 0),
		(drawing, 1444, 0, 2048, 0, 0),
		(drawing, 1445, 0, 2048, 0, 0),
		(drawing, 1446, 0, 2048, 0, 0),
		(drawing, 1447, 0, 2048, 0, 0),
		(drawing, 1448, 0, 2048, 0, 0),
		(drawing, 1449, 0, 2048, 0, 0),
		(drawing, 1450, 0, 2048, 0, 0),
		(drawing, 1451, 0, 2048, 0, 0),
		(drawing, 1452, 0, 2048, 0, 0),
		(drawing, 1453, 0, 2048, 0, 0),
		(drawing, 1454, 0, 2048, 0, 0),
		(drawing, 1455, 0, 2048, 0, 0),
		(drawing, 1456, 0, 2048, 0, 0),
		(drawing, 1457, 0, 2048, 0, 0),
		(drawing, 1458, 0, 2048, 0, 0),
		(drawing, 1459, 0, 2048, 0, 0),
		(drawing, 1460, 0, 2048, 0, 0),
		(drawing, 1461, 0, 2048, 0, 0),
		(drawing, 1462, 0, 2048, 0, 0),
		(drawing, 1463, 0, 2048, 0, 0),
		(drawing, 1464, 0, 2048, 0, 0),
		(drawing, 1465, 0, 2048, 0, 0),
		(drawing, 1466, 0, 2048, 0, 0),
		(drawing, 1467, 0, 2048, 0, 0),
		(drawing, 1468, 0, 2048, 0, 0),
		(drawing, 1469, 0, 2048, 0, 0),
		(drawing, 1470, 0, 2048, 0, 0),
		(drawing, 1471, 0, 2048, 0, 0),
		(drawing, 1472, 0, 2048, 0, 0),
		(drawing, 1473, 0, 2048, 0, 0),
		(drawing, 1474, 0, 2048, 0, 0),
		(drawing, 1475, 0, 2048, 0, 0),
		(drawing, 1476, 0, 2048, 0, 0),
		(drawing, 1477, 0, 2048, 0, 0),
		(drawing, 1478, 0, 2048, 0, 0),
		(drawing, 1479, 0, 2048, 0, 0),
		(drawing, 1480, 0, 2048, 0, 0),
		(drawing, 1481, 0, 2048, 0, 0),
		(drawing, 1482, 0, 2048, 0, 0),
		(drawing, 1483, 0, 2048, 0, 0),
		(drawing, 1484, 0, 2048, 0, 0),
		(drawing, 1485, 0, 2048, 0, 0),
		(drawing, 1486, 0, 2048, 0, 0),
		(drawing, 1487, 0, 2048, 0, 0),
		(drawing, 1488, 0, 2048, 0, 0),
		(drawing, 1489, 0, 2048, 0, 0),
		(drawing, 1490, 0, 2048, 0, 0),
		(drawing, 1491, 0, 2048, 0, 0),
		(drawing, 1492, 0, 2048, 0, 0),
		(drawing, 1493, 0, 2048, 0, 0),
		(drawing, 1494, 0, 2048, 0, 0),
		(drawing, 1495, 0, 2048, 0, 0),
		(drawing, 1496, 0, 2048, 0, 0),
		(drawing, 1497, 0, 2048, 0, 0),
		(drawing, 1498, 0, 2048, 0, 0),
		(drawing, 1499, 0, 2048, 0, 0),
		(drawing, 1500, 0, 2048, 0, 0),
		(drawing, 1501, 0, 2048, 0, 0),
		(drawing, 1502, 0, 2048, 0, 0),
		(drawing, 1503, 0, 2048, 0, 0),
		(drawing, 1504, 0, 2048, 0, 0),
		(drawing, 1505, 0, 2048, 0, 0),
		(drawing, 1506, 0, 2048, 0, 0),
		(drawing, 1507, 0, 2048, 0, 0),
		(drawing, 1508, 0, 2048, 0, 0),
		(drawing, 1509, 0, 2048, 0, 0),
		(drawing, 1510, 0, 2048, 0, 0),
		(drawing, 1511, 0, 2048, 0, 0),
		(drawing, 1512, 0, 2048, 0, 0),
		(drawing, 1513, 0, 2048, 0, 0),
		(drawing, 1514, 0, 2048, 0, 0),
		(drawing, 1515, 0, 2048, 0, 0),
		(drawing, 1516, 0, 2048, 0, 0),
		(drawing, 1517, 0, 2048, 0, 0),
		(drawing, 1518, 0, 2048, 0, 0),
		(drawing, 1519, 0, 2048, 0, 0),
		(drawing, 1520, 0, 2048, 0, 0),
		(drawing, 1521, 0, 2048, 0, 0),
		(drawing, 1522, 0, 2048, 0, 0),
		(drawing, 1523, 0, 2048, 0, 0),
		(drawing, 1524, 0, 2048, 0, 0),
		(drawing, 1525, 0, 2048, 0, 0),
		(drawing, 1526, 0, 2048, 0, 0),
		(drawing, 1527, 0, 2048, 0, 0),
		(drawing, 1528, 0, 2048, 0, 0),
		(drawing, 1529, 0, 2048, 0, 0),
		(drawing, 1530, 0, 2048, 0, 0),
		(drawing, 1531, 0, 2048, 0, 0),
		(drawing, 1532, 0, 2048, 0, 0),
		(drawing, 1533, 0, 2048, 0, 0),
		(drawing, 1534, 0, 2048, 0, 0),
		(drawing, 1535, 0, 2048, 0, 0),
		(drawing, 1536, 0, 2048, 0, 0),
		(drawing, 1537, 0, 2048, 0, 0),
		(drawing, 1538, 0, 2048, 0, 0),
		(drawing, 1539, 0, 2048, 0, 0),
		(drawing, 1540, 0, 2048, 0, 0),
		(drawing, 1541, 0, 2048, 0, 0),
		(drawing, 1542, 0, 2048, 0, 0),
		(drawing, 1543, 0, 2048, 0, 0),
		(drawing, 1544, 0, 2048, 0, 0),
		(drawing, 1545, 0, 2048, 0, 0),
		(drawing, 1546, 0, 2048, 0, 0),
		(drawing, 1547, 0, 2048, 0, 0),
		(drawing, 1548, 0, 2048, 0, 0),
		(drawing, 1549, 0, 2048, 0, 0),
		(drawing, 1550, 0, 2048, 0, 0),
		(drawing, 1551, 0, 2048, 0, 0),
		(drawing, 1552, 0, 2048, 0, 0),
		(drawing, 1553, 0, 2048, 0, 0),
		(drawing, 1554, 0, 2048, 0, 0),
		(drawing, 1555, 0, 2048, 0, 0),
		(drawing, 1556, 0, 2048, 0, 0),
		(drawing, 1557, 0, 2048, 0, 0),
		(drawing, 1558, 0, 2048, 0, 0),
		(drawing, 1559, 0, 2048, 0, 0),
		(drawing, 1560, 0, 2048, 0, 0),
		(drawing, 1561, 0, 2048, 0, 0),
		(drawing, 1562, 0, 2048, 0, 0),
		(drawing, 1563, 0, 2048, 0, 0),
		(drawing, 1564, 0, 2048, 0, 0),
		(drawing, 1565, 0, 2048, 0, 0),
		(drawing, 1566, 0, 2048, 0, 0),
		(drawing, 1567, 0, 2048, 0, 0),
		(drawing, 1568, 0, 2048, 0, 0),
		(drawing, 1569, 0, 2048, 0, 0),
		(drawing, 1570, 0, 2048, 0, 0),
		(drawing, 1571, 0, 2048, 0, 0),
		(drawing, 1572, 0, 2048, 0, 0),
		(drawing, 1573, 0, 2048, 0, 0),
		(drawing, 1574, 0, 2048, 0, 0),
		(drawing, 1575, 0, 2048, 0, 0),
		(drawing, 1576, 0, 2048, 0, 0),
		(drawing, 1577, 0, 2048, 0, 0),
		(drawing, 1578, 0, 2048, 0, 0),
		(drawing, 1579, 0, 2048, 0, 0),
		(drawing, 1580, 0, 2048, 0, 0),
		(drawing, 1581, 0, 2048, 0, 0),
		(drawing, 1582, 0, 2048, 0, 0),
		(drawing, 1583, 0, 2048, 0, 0),
		(drawing, 1584, 0, 2048, 0, 0),
		(drawing, 1585, 0, 2048, 0, 0),
		(drawing, 1586, 0, 2048, 0, 0),
		(drawing, 1587, 0, 2048, 0, 0),
		(drawing, 1588, 0, 2048, 0, 0),
		(drawing, 1589, 0, 2048, 0, 0),
		(drawing, 1590, 0, 2048, 0, 0),
		(drawing, 1591, 0, 2048, 0, 0),
		(drawing, 1592, 0, 2048, 0, 0),
		(drawing, 1593, 0, 2048, 0, 0),
		(drawing, 1594, 0, 2048, 0, 0),
		(drawing, 1595, 0, 2048, 0, 0),
		(drawing, 1596, 0, 2048, 0, 0),
		(drawing, 1597, 0, 2048, 0, 0),
		(drawing, 1598, 0, 2048, 0, 0),
		(drawing, 1599, 0, 2048, 0, 0),
		(drawing, 1600, 0, 2048, 0, 0),
		(drawing, 1601, 0, 2048, 0, 0),
		(drawing, 1602, 0, 2048, 0, 0),
		(drawing, 1603, 0, 2048, 0, 0),
		(drawing, 1604, 0, 2048, 0, 0),
		(drawing, 1605, 0, 2048, 0, 0),
		(drawing, 1606, 0, 2048, 0, 0),
		(drawing, 1607, 0, 2048, 0, 0),
		(drawing, 1608, 0, 2048, 0, 0),
		(drawing, 1609, 0, 2048, 0, 0),
		(drawing, 1610, 0, 2048, 0, 0),
		(drawing, 1611, 0, 2048, 0, 0),
		(drawing, 1612, 0, 2048, 0, 0),
		(drawing, 1613, 0, 2048, 0, 0),
		(drawing, 1614, 0, 2048, 0, 0),
		(drawing, 1615, 0, 2048, 0, 0),
		(drawing, 1616, 0, 2048, 0, 0),
		(drawing, 1617, 0, 2048, 0, 0),
		(drawing, 1618, 0, 2048, 0, 0),
		(drawing, 1619, 0, 2048, 0, 0),
		(drawing, 1620, 0, 2048, 0, 0),
		(drawing, 1621, 0, 2048, 0, 0),
		(drawing, 1622, 0, 2048, 0, 0),
		(drawing, 1623, 0, 2048, 0, 0),
		(drawing, 1624, 0, 2048, 0, 0),
		(drawing, 1625, 0, 2048, 0, 0),
		(drawing, 1626, 0, 2048, 0, 0),
		(drawing, 1627, 0, 2048, 0, 0),
		(drawing, 1628, 0, 2048, 0, 0),
		(drawing, 1629, 0, 2048, 0, 0),
		(drawing, 1630, 0, 2048, 0, 0),
		(drawing, 1631, 0, 2048, 0, 0),
		(drawing, 1632, 0, 2048, 0, 0),
		(drawing, 1633, 0, 2048, 0, 0),
		(drawing, 1634, 0, 2048, 0, 0),
		(drawing, 1635, 0, 2048, 0, 0),
		(drawing, 1636, 0, 2048, 0, 0),
		(drawing, 1637, 0, 2048, 0, 0),
		(drawing, 1638, 0, 2048, 0, 0),
		(drawing, 1639, 0, 2048, 0, 0),
		(drawing, 1640, 0, 2048, 0, 0),
		(drawing, 1641, 0, 2048, 0, 0),
		(drawing, 1642, 0, 2048, 0, 0),
		(drawing, 1643, 0, 2048, 0, 0),
		(drawing, 1644, 0, 2048, 0, 0),
		(drawing, 1645, 0, 2048, 0, 0),
		(drawing, 1646, 0, 2048, 0, 0),
		(drawing, 1647, 0, 2048, 0, 0),
		(drawing, 1648, 0, 2048, 0, 0),
		(drawing, 1649, 0, 2048, 0, 0),
		(drawing, 1650, 0, 2048, 0, 0),
		(drawing, 1651, 0, 2048, 0, 0),
		(drawing, 1652, 0, 2048, 0, 0),
		(drawing, 1653, 0, 2048, 0, 0),
		(drawing, 1654, 0, 2048, 0, 0),
		(drawing, 1655, 0, 2048, 0, 0),
		(drawing, 1656, 0, 2048, 0, 0),
		(drawing, 1657, 0, 2048, 0, 0),
		(drawing, 1658, 0, 2048, 0, 0),
		(drawing, 1659, 0, 2048, 0, 0),
		(drawing, 1660, 0, 2048, 0, 0),
		(drawing, 1661, 0, 2048, 0, 0),
		(drawing, 1662, 0, 2048, 0, 0),
		(drawing, 1663, 0, 2048, 0, 0),
		(drawing, 1664, 0, 2048, 0, 0),
		(drawing, 1665, 0, 2048, 0, 0),
		(drawing, 1666, 0, 2048, 0, 0),
		(drawing, 1667, 0, 2048, 0, 0),
		(drawing, 1668, 0, 2048, 0, 0),
		(drawing, 1669, 0, 2048, 0, 0),
		(drawing, 1670, 0, 2048, 0, 0),
		(drawing, 1671, 0, 2048, 0, 0),
		(drawing, 1672, 0, 2048, 0, 0),
		(drawing, 1673, 0, 2048, 0, 0),
		(drawing, 1674, 0, 2048, 0, 0),
		(drawing, 1675, 0, 2048, 0, 0),
		(drawing, 1676, 0, 2048, 0, 0),
		(drawing, 1677, 0, 2048, 0, 0),
		(drawing, 1678, 0, 2048, 0, 0),
		(drawing, 1679, 0, 2048, 0, 0),
		(drawing, 1680, 0, 2048, 0, 0),
		(drawing, 1681, 0, 2048, 0, 0),
		(drawing, 1682, 0, 2048, 0, 0),
		(drawing, 1683, 0, 2048, 0, 0),
		(drawing, 1684, 0, 2048, 0, 0),
		(drawing, 1685, 0, 2048, 0, 0),
		(drawing, 1686, 0, 2048, 0, 0),
		(drawing, 1687, 0, 2048, 0, 0),
		(drawing, 1688, 0, 2048, 0, 0),
		(drawing, 1689, 0, 2048, 0, 0),
		(drawing, 1690, 0, 2048, 0, 0),
		(drawing, 1691, 0, 2048, 0, 0),
		(drawing, 1692, 0, 2048, 0, 0),
		(drawing, 1693, 0, 2048, 0, 0),
		(drawing, 1694, 0, 2048, 0, 0),
		(drawing, 1695, 0, 2048, 0, 0),
		(drawing, 1696, 0, 2048, 0, 0),
		(drawing, 1697, 0, 2048, 0, 0),
		(drawing, 1698, 0, 2048, 0, 0),
		(drawing, 1699, 0, 2048, 0, 0),
		(drawing, 1700, 0, 2048, 0, 0),
		(drawing, 1701, 0, 2048, 0, 0),
		(drawing, 1702, 0, 2048, 0, 0),
		(drawing, 1703, 0, 2048, 0, 0),
		(drawing, 1704, 0, 2048, 0, 0),
		(drawing, 1705, 0, 2048, 0, 0),
		(drawing, 1706, 0, 2048, 0, 0),
		(drawing, 1707, 0, 2048, 0, 0),
		(drawing, 1708, 0, 2048, 0, 0),
		(drawing, 1709, 0, 2048, 0, 0),
		(drawing, 1710, 0, 2048, 0, 0),
		(drawing, 1711, 0, 2048, 0, 0),
		(drawing, 1712, 0, 2048, 0, 0),
		(drawing, 1713, 0, 2048, 0, 0),
		(drawing, 1714, 0, 2048, 0, 0),
		(drawing, 1715, 0, 2048, 0, 0),
		(drawing, 1716, 0, 2048, 0, 0),
		(drawing, 1717, 0, 2048, 0, 0),
		(drawing, 1718, 0, 2048, 0, 0),
		(drawing, 1719, 0, 2048, 0, 0),
		(drawing, 1720, 0, 2048, 0, 0),
		(drawing, 1721, 0, 2048, 0, 0),
		(drawing, 1722, 0, 2048, 0, 0),
		(drawing, 1723, 0, 2048, 0, 0),
		(drawing, 1724, 0, 2048, 0, 0),
		(drawing, 1725, 0, 2048, 0, 0),
		(drawing, 1726, 0, 2048, 0, 0),
		(drawing, 1727, 0, 2048, 0, 0),
		(drawing, 1728, 0, 2048, 0, 0),
		(drawing, 1729, 0, 2048, 0, 0),
		(drawing, 1730, 0, 2048, 0, 0),
		(drawing, 1731, 0, 2048, 0, 0),
		(drawing, 1732, 0, 2048, 0, 0),
		(drawing, 1733, 0, 2048, 0, 0),
		(drawing, 1734, 0, 2048, 0, 0),
		(drawing, 1735, 0, 2048, 0, 0),
		(drawing, 1736, 0, 2048, 0, 0),
		(drawing, 1737, 0, 2048, 0, 0),
		(drawing, 1738, 0, 2048, 0, 0),
		(drawing, 1739, 0, 2048, 0, 0),
		(drawing, 1740, 0, 2048, 0, 0),
		(drawing, 1741, 0, 2048, 0, 0),
		(drawing, 1742, 0, 2048, 0, 0),
		(drawing, 1743, 0, 2048, 0, 0),
		(drawing, 1744, 0, 2048, 0, 0),
		(drawing, 1745, 0, 2048, 0, 0),
		(drawing, 1746, 0, 2048, 0, 0),
		(drawing, 1747, 0, 2048, 0, 0),
		(drawing, 1748, 0, 2048, 0, 0),
		(drawing, 1749, 0, 2048, 0, 0),
		(drawing, 1750, 0, 2048, 0, 0),
		(drawing, 1751, 0, 2048, 0, 0),
		(drawing, 1752, 0, 2048, 0, 0),
		(drawing, 1753, 0, 2048, 0, 0),
		(drawing, 1754, 0, 2048, 0, 0),
		(drawing, 1755, 0, 2048, 0, 0),
		(drawing, 1756, 0, 2048, 0, 0),
		(drawing, 1757, 0, 2048, 0, 0),
		(drawing, 1758, 0, 2048, 0, 0),
		(drawing, 1759, 0, 2048, 0, 0),
		(drawing, 1760, 0, 2048, 0, 0),
		(drawing, 1761, 0, 2048, 0, 0),
		(drawing, 1762, 0, 2048, 0, 0),
		(drawing, 1763, 0, 2048, 0, 0),
		(drawing, 1764, 0, 2048, 0, 0),
		(drawing, 1765, 0, 2048, 0, 0),
		(drawing, 1766, 0, 2048, 0, 0),
		(drawing, 1767, 0, 2048, 0, 0),
		(drawing, 1768, 0, 2048, 0, 0),
		(drawing, 1769, 0, 2048, 0, 0),
		(drawing, 1770, 0, 2048, 0, 0),
		(drawing, 1771, 0, 2048, 0, 0),
		(drawing, 1772, 0, 2048, 0, 0),
		(drawing, 1773, 0, 2048, 0, 0),
		(drawing, 1774, 0, 2048, 0, 0),
		(drawing, 1775, 0, 2048, 0, 0),
		(drawing, 1776, 0, 2048, 0, 0),
		(drawing, 1777, 0, 2048, 0, 0),
		(drawing, 1778, 0, 2048, 0, 0),
		(drawing, 1779, 0, 2048, 0, 0),
		(drawing, 1780, 0, 2048, 0, 0),
		(drawing, 1781, 0, 2048, 0, 0),
		(drawing, 1782, 0, 2048, 0, 0),
		(drawing, 1783, 0, 2048, 0, 0),
		(drawing, 1784, 0, 2048, 0, 0),
		(drawing, 1785, 0, 2048, 0, 0),
		(drawing, 1786, 0, 2048, 0, 0),
		(drawing, 1787, 0, 2048, 0, 0),
		(drawing, 1788, 0, 2048, 0, 0),
		(drawing, 1789, 0, 2048, 0, 0),
		(drawing, 1790, 0, 2048, 0, 0),
		(drawing, 1791, 0, 2048, 0, 0),
		(drawing, 1792, 0, 2048, 0, 0),
		(drawing, 1793, 0, 2048, 0, 0),
		(drawing, 1794, 0, 2048, 0, 0),
		(drawing, 1795, 0, 2048, 0, 0),
		(drawing, 1796, 0, 2048, 0, 0),
		(drawing, 1797, 0, 2048, 0, 0),
		(drawing, 1798, 0, 2048, 0, 0),
		(drawing, 1799, 0, 2048, 0, 0),
		(drawing, 1800, 0, 2048, 0, 0),
		(drawing, 1801, 0, 2048, 0, 0),
		(drawing, 1802, 0, 2048, 0, 0),
		(drawing, 1803, 0, 2048, 0, 0),
		(drawing, 1804, 0, 2048, 0, 0),
		(drawing, 1805, 0, 2048, 0, 0),
		(drawing, 1806, 0, 2048, 0, 0),
		(drawing, 1807, 0, 2048, 0, 0),
		(drawing, 1808, 0, 2048, 0, 0),
		(drawing, 1809, 0, 2048, 0, 0),
		(drawing, 1810, 0, 2048, 0, 0),
		(drawing, 1811, 0, 2048, 0, 0),
		(drawing, 1812, 0, 2048, 0, 0),
		(drawing, 1813, 0, 2048, 0, 0),
		(drawing, 1814, 0, 2048, 0, 0),
		(drawing, 1815, 0, 2048, 0, 0),
		(drawing, 1816, 0, 2048, 0, 0),
		(drawing, 1817, 0, 2048, 0, 0),
		(drawing, 1818, 0, 2048, 0, 0),
		(drawing, 1819, 0, 2048, 0, 0),
		(drawing, 1820, 0, 2048, 0, 0),
		(drawing, 1821, 0, 2048, 0, 0),
		(drawing, 1822, 0, 2048, 0, 0),
		(drawing, 1823, 0, 2048, 0, 0),
		(drawing, 1824, 0, 2048, 0, 0),
		(drawing, 1825, 0, 2048, 0, 0),
		(drawing, 1826, 0, 2048, 0, 0),
		(drawing, 1827, 0, 2048, 0, 0),
		(drawing, 1828, 0, 2048, 0, 0),
		(drawing, 1829, 0, 2048, 0, 0),
		(drawing, 1830, 0, 2048, 0, 0),
		(drawing, 1831, 0, 2048, 0, 0),
		(drawing, 1832, 0, 2048, 0, 0),
		(drawing, 1833, 0, 2048, 0, 0),
		(drawing, 1834, 0, 2048, 0, 0),
		(drawing, 1835, 0, 2048, 0, 0),
		(drawing, 1836, 0, 2048, 0, 0),
		(drawing, 1837, 0, 2048, 0, 0),
		(drawing, 1838, 0, 2048, 0, 0),
		(drawing, 1839, 0, 2048, 0, 0),
		(drawing, 1840, 0, 2048, 0, 0),
		(drawing, 1841, 0, 2048, 0, 0),
		(drawing, 1842, 0, 2048, 0, 0),
		(drawing, 1843, 0, 2048, 0, 0),
		(drawing, 1844, 0, 2048, 0, 0),
		(drawing, 1845, 0, 2048, 0, 0),
		(drawing, 1846, 0, 2048, 0, 0),
		(drawing, 1847, 0, 2048, 0, 0),
		(drawing, 1848, 0, 2048, 0, 0),
		(drawing, 1849, 0, 2048, 0, 0),
		(drawing, 1850, 0, 2048, 0, 0),
		(drawing, 1851, 0, 2048, 0, 0),
		(drawing, 1852, 0, 2048, 0, 0),
		(drawing, 1853, 0, 2048, 0, 0),
		(drawing, 1854, 0, 2048, 0, 0),
		(drawing, 1855, 0, 2048, 0, 0),
		(drawing, 1856, 0, 2048, 0, 0),
		(drawing, 1857, 0, 2048, 0, 0),
		(drawing, 1858, 0, 2048, 0, 0),
		(drawing, 1859, 0, 2048, 0, 0),
		(drawing, 1860, 0, 2048, 0, 0),
		(drawing, 1861, 0, 2048, 0, 0),
		(drawing, 1862, 0, 2048, 0, 0),
		(drawing, 1863, 0, 2048, 0, 0),
		(drawing, 1864, 0, 2048, 0, 0),
		(drawing, 1865, 0, 2048, 0, 0),
		(drawing, 1866, 0, 2048, 0, 0),
		(drawing, 1867, 0, 2048, 0, 0),
		(drawing, 1868, 0, 2048, 0, 0),
		(drawing, 1869, 0, 2048, 0, 0),
		(drawing, 1870, 0, 2048, 0, 0),
		(drawing, 1871, 0, 2048, 0, 0),
		(drawing, 1872, 0, 2048, 0, 0),
		(drawing, 1873, 0, 2048, 0, 0),
		(drawing, 1874, 0, 2048, 0, 0),
		(drawing, 1875, 0, 2048, 0, 0),
		(drawing, 1876, 0, 2048, 0, 0),
		(drawing, 1877, 0, 2048, 0, 0),
		(drawing, 1878, 0, 2048, 0, 0),
		(drawing, 1879, 0, 2048, 0, 0),
		(drawing, 1880, 0, 2048, 0, 0),
		(drawing, 1881, 0, 2048, 0, 0),
		(drawing, 1882, 0, 2048, 0, 0),
		(drawing, 1883, 0, 2048, 0, 0),
		(drawing, 1884, 0, 2048, 0, 0),
		(drawing, 1885, 0, 2048, 0, 0),
		(drawing, 1886, 0, 2048, 0, 0),
		(drawing, 1887, 0, 2048, 0, 0),
		(drawing, 1888, 0, 2048, 0, 0),
		(drawing, 1889, 0, 2048, 0, 0),
		(drawing, 1890, 0, 2048, 0, 0),
		(drawing, 1891, 0, 2048, 0, 0),
		(drawing, 1892, 0, 2048, 0, 0),
		(drawing, 1893, 0, 2048, 0, 0),
		(drawing, 1894, 0, 2048, 0, 0),
		(drawing, 1895, 0, 2048, 0, 0),
		(drawing, 1896, 0, 2048, 0, 0),
		(drawing, 1897, 0, 2048, 0, 0),
		(drawing, 1898, 0, 2048, 0, 0),
		(drawing, 1899, 0, 2048, 0, 0),
		(drawing, 1900, 0, 2048, 0, 0),
		(drawing, 1901, 0, 2048, 0, 0),
		(drawing, 1902, 0, 2048, 0, 0),
		(drawing, 1903, 0, 2048, 0, 0),
		(drawing, 1904, 0, 2048, 0, 0),
		(drawing, 1905, 0, 2048, 0, 0),
		(drawing, 1906, 0, 2048, 0, 0),
		(drawing, 1907, 0, 2048, 0, 0),
		(drawing, 1908, 0, 2048, 0, 0),
		(drawing, 1909, 0, 2048, 0, 0),
		(drawing, 1910, 0, 2048, 0, 0),
		(drawing, 1911, 0, 2048, 0, 0),
		(drawing, 1912, 0, 2048, 0, 0),
		(drawing, 1913, 0, 2048, 0, 0),
		(drawing, 1914, 0, 2048, 0, 0),
		(drawing, 1915, 0, 2048, 0, 0),
		(drawing, 1916, 0, 2048, 0, 0),
		(drawing, 1917, 0, 2048, 0, 0),
		(drawing, 1918, 0, 2048, 0, 0),
		(drawing, 1919, 0, 2048, 0, 0),
		(drawing, 1920, 0, 2048, 0, 0),
		(drawing, 1921, 0, 2048, 0, 0),
		(drawing, 1922, 0, 2048, 0, 0),
		(drawing, 1923, 0, 2048, 0, 0),
		(drawing, 1924, 0, 2048, 0, 0),
		(drawing, 1925, 0, 2048, 0, 0),
		(drawing, 1926, 0, 2048, 0, 0),
		(drawing, 1927, 0, 2048, 0, 0),
		(drawing, 1928, 0, 2048, 0, 0),
		(drawing, 1929, 0, 2048, 0, 0),
		(drawing, 1930, 0, 2048, 0, 0),
		(drawing, 1931, 0, 2048, 0, 0),
		(drawing, 1932, 0, 2048, 0, 0),
		(drawing, 1933, 0, 2048, 0, 0),
		(drawing, 1934, 0, 2048, 0, 0),
		(drawing, 1935, 0, 2048, 0, 0),
		(drawing, 1936, 0, 2048, 0, 0),
		(drawing, 1937, 0, 2048, 0, 0),
		(drawing, 1938, 0, 2048, 0, 0),
		(drawing, 1939, 0, 2048, 0, 0),
		(drawing, 1940, 0, 2048, 0, 0),
		(drawing, 1941, 0, 2048, 0, 0),
		(drawing, 1942, 0, 2048, 0, 0),
		(drawing, 1943, 0, 2048, 0, 0),
		(drawing, 1944, 0, 2048, 0, 0),
		(drawing, 1945, 0, 2048, 0, 0),
		(drawing, 1946, 0, 2048, 0, 0),
		(drawing, 1947, 0, 2048, 0, 0),
		(drawing, 1948, 0, 2048, 0, 0),
		(drawing, 1949, 0, 2048, 0, 0),
		(drawing, 1950, 0, 2048, 0, 0),
		(drawing, 1951, 0, 2048, 0, 0),
		(drawing, 1952, 0, 2048, 0, 0),
		(drawing, 1953, 0, 2048, 0, 0),
		(drawing, 1954, 0, 2048, 0, 0),
		(drawing, 1955, 0, 2048, 0, 0),
		(drawing, 1956, 0, 2048, 0, 0),
		(drawing, 1957, 0, 2048, 0, 0),
		(drawing, 1958, 0, 2048, 0, 0),
		(drawing, 1959, 0, 2048, 0, 0),
		(drawing, 1960, 0, 2048, 0, 0),
		(drawing, 1961, 0, 2048, 0, 0),
		(drawing, 1962, 0, 2048, 0, 0),
		(drawing, 1963, 0, 2048, 0, 0),
		(drawing, 1964, 0, 2048, 0, 0),
		(drawing, 1965, 0, 2048, 0, 0),
		(drawing, 1966, 0, 2048, 0, 0),
		(drawing, 1967, 0, 2048, 0, 0),
		(drawing, 1968, 0, 2048, 0, 0),
		(drawing, 1969, 0, 2048, 0, 0),
		(drawing, 1970, 0, 2048, 0, 0),
		(drawing, 1971, 0, 2048, 0, 0),
		(drawing, 1972, 0, 2048, 0, 0),
		(drawing, 1973, 0, 2048, 0, 0),
		(drawing, 1974, 0, 2048, 0, 0),
		(drawing, 1975, 0, 2048, 0, 0),
		(drawing, 1976, 0, 2048, 0, 0),
		(drawing, 1977, 0, 2048, 0, 0),
		(drawing, 1978, 0, 2048, 0, 0),
		(drawing, 1979, 0, 2048, 0, 0),
		(drawing, 1980, 0, 2048, 0, 0),
		(drawing, 1981, 0, 2048, 0, 0),
		(drawing, 1982, 0, 2048, 0, 0),
		(drawing, 1983, 0, 2048, 0, 0),
		(drawing, 1984, 0, 2048, 0, 0),
		(drawing, 1985, 0, 2048, 0, 0),
		(drawing, 1986, 0, 2048, 0, 0),
		(drawing, 1987, 0, 2048, 0, 0),
		(drawing, 1988, 0, 2048, 0, 0),
		(drawing, 1989, 0, 2048, 0, 0),
		(drawing, 1990, 0, 2048, 0, 0),
		(drawing, 1991, 0, 2048, 0, 0),
		(drawing, 1992, 0, 2048, 0, 0),
		(drawing, 1993, 0, 2048, 0, 0),
		(drawing, 1994, 0, 2048, 0, 0),
		(drawing, 1995, 0, 2048, 0, 0),
		(drawing, 1996, 0, 2048, 0, 0),
		(drawing, 1997, 0, 2048, 0, 0),
		(drawing, 1998, 0, 2048, 0, 0),
		(drawing, 1999, 0, 2048, 0, 0),
		(drawing, 2000, 0, 2048, 0, 0),
		(drawing, 2001, 0, 2048, 0, 0),
		(drawing, 2002, 0, 2048, 0, 0),
		(drawing, 2003, 0, 2048, 0, 0),
		(drawing, 2004, 0, 2048, 0, 0),
		(drawing, 2005, 0, 2048, 0, 0),
		(drawing, 2006, 0, 2048, 0, 0),
		(drawing, 2007, 0, 2048, 0, 0),
		(drawing, 2008, 0, 2048, 0, 0),
		(drawing, 2009, 0, 2048, 0, 0),
		(drawing, 2010, 0, 2048, 0, 0),
		(drawing, 2011, 0, 2048, 0, 0),
		(drawing, 2012, 0, 2048, 0, 0),
		(drawing, 2013, 0, 2048, 0, 0),
		(drawing, 2014, 0, 2048, 0, 0),
		(drawing, 2015, 0, 2048, 0, 0),
		(drawing, 2016, 0, 2048, 0, 0),
		(drawing, 2017, 0, 2048, 0, 0),
		(drawing, 2018, 0, 2048, 0, 0),
		(drawing, 2019, 0, 2048, 0, 0),
		(drawing, 2020, 0, 2048, 0, 0),
		(drawing, 2021, 0, 2048, 0, 0),
		(drawing, 2022, 0, 2048, 0, 0),
		(drawing, 2023, 0, 2048, 0, 0),
		(drawing, 2024, 0, 2048, 0, 0),
		(drawing, 2025, 0, 2048, 0, 0),
		(drawing, 2026, 0, 2048, 0, 0),
		(drawing, 2027, 0, 2048, 0, 0),
		(drawing, 2028, 0, 2048, 0, 0),
		(drawing, 2029, 0, 2048, 0, 0),
		(drawing, 2030, 0, 2048, 0, 0),
		(drawing, 2031, 0, 2048, 0, 0),
		(drawing, 2032, 0, 2048, 0, 0),
		(drawing, 2033, 0, 2048, 0, 0),
		(drawing, 2034, 0, 2048, 0, 0),
		(drawing, 2035, 0, 2048, 0, 0),
		(drawing, 2036, 0, 2048, 0, 0),
		(drawing, 2037, 0, 2048, 0, 0),
		(drawing, 2038, 0, 2048, 0, 0),
		(drawing, 2039, 0, 2048, 0, 0),
		(drawing, 2040, 0, 2048, 0, 0),
		(drawing, 2041, 0, 2048, 0, 0),
		(drawing, 2042, 0, 2048, 0, 0),
		(drawing, 2043, 0, 2048, 0, 0),
		(drawing, 2044, 0, 2048, 0, 0),
		(drawing, 2045, 0, 2048, 0, 0),
		(drawing, 2046, 0, 2048, 0, 0),
		(drawing, 2047, 0, 2048, 0, 0),
		(done, 2048, 0, 2048, 0, 0)
	);
END PACKAGE ex1_data_pak;
