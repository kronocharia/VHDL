
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE WORK.pix_cache_pak.ALL;
USE WORK.pix_tb_pak.ALL;

PACKAGE ex4_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        rst,wen_all,pw: INTEGER;
        pixop:  pixop_tb_t;
        pixnum: INTEGER;
        is_same: INTEGER;
        store: pixop_tb_vec(0 TO 15);
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(
--                 INPUTS              ||           OUTPUTS
--  rst    wen_all  pw   pixop pixnum      is_same   store

	(1,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     0,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     11,     0, "W:::::W:::::::::"),
	(0,     0,     1,     '*',     11,     0, "W:::::W::::W::::"),
	(0,     0,     0,     ':',     7,     0, "W:::::W::::B::::"),
	(0,     0,     0,     ':',     2,     0, "W:::::W::::B::::"),
	(0,     0,     0,     ':',     5,     0, "W:::::W::::B::::"),
	(0,     0,     1,     'B',     14,     0, "W:::::W::::B::::"),
	(0,     0,     0,     'B',     12,     0, "W:::::W::::B::B:"),
	(0,     0,     0,     ':',     9,     0, "W:::::W::::B::B:"),
	(0,     0,     1,     'B',     8,     0, "W:::::W::::B::B:"),
	(0,     0,     1,     ':',     0,     0, "W:::::W:B::B::B:"),
	(0,     1,     0,     ':',     3,     0, "W:::::W:B::B::B:"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     0, ":::::::W::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::::BW::::::::"),
	(0,     0,     1,     'B',     9,     0, "::::::BW::::::::"),
	(0,     0,     0,     'B',     12,     0, "::::::BW:B::::::"),
	(0,     0,     1,     'W',     7,     0, "::::::BW:B::::::"),
	(0,     0,     1,     'B',     14,     0, "::::::BW:B::::::"),
	(0,     0,     0,     '*',     10,     0, "::::::BW:B::::B:"),
	(0,     0,     0,     ':',     9,     0, "::::::BW:B::::B:"),
	(0,     0,     1,     'W',     12,     0, "::::::BW:B::::B:"),
	(0,     0,     0,     '*',     2,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     'B',     8,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     ':',     11,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     ':',     9,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     'B',     14,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     '*',     1,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     'B',     10,     0, "::::::BW:B::W:B:"),
	(1,     0,     0,     'B',     2,     0, "::::::BW:B::W:B:"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     13,     0, ":::::B::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::::B:::::::B::"),
	(0,     0,     1,     'B',     10,     0, ":::::B:::::::B::"),
	(0,     0,     1,     'B',     1,     0, ":::::B::::B::B::"),
	(0,     0,     0,     'B',     8,     0, ":B:::B::::B::B::"),
	(0,     1,     0,     'B',     6,     0, ":B:::B::::B::B::"),
	(0,     1,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     0, "::B:::::::::::::"),
	(0,     0,     0,     'B',     9,     0, "::B:::::::::::::"),
	(0,     0,     1,     'W',     11,     0, "::B:::::::::::::"),
	(0,     0,     1,     'W',     0,     0, "::B::::::::W::::"),
	(0,     0,     1,     ':',     9,     0, "W:B::::::::W::::"),
	(0,     0,     1,     'W',     14,     0, "W:B::::::::W::::"),
	(0,     0,     1,     '*',     9,     0, "W:B::::::::W::W:"),
	(0,     0,     0,     ':',     11,     0, "W:B::::::*:W::W:"),
	(0,     0,     1,     'B',     6,     0, "W:B::::::*:W::W:"),
	(0,     0,     0,     'B',     9,     0, "W:B:::B::*:W::W:"),
	(0,     0,     1,     'W',     11,     0, "W:B:::B::*:W::W:"),
	(0,     0,     1,     'B',     13,     0, "W:B:::B::*:W::W:"),
	(0,     0,     0,     'B',     7,     0, "W:B:::B::*:W:BW:"),
	(0,     0,     0,     '*',     7,     0, "W:B:::B::*:W:BW:"),
	(0,     0,     1,     'B',     1,     0, "W:B:::B::*:W:BW:"),
	(0,     0,     0,     'B',     9,     0, "WBB:::B::*:W:BW:"),
	(0,     0,     1,     '*',     2,     0, "WBB:::B::*:W:BW:"),
	(0,     0,     0,     'W',     7,     0, "WBW:::B::*:W:BW:"),
	(0,     0,     0,     ':',     2,     0, "WBW:::B::*:W:BW:"),
	(0,     0,     0,     ':',     10,     0, "WBW:::B::*:W:BW:"),
	(0,     0,     1,     '*',     9,     0, "WBW:::B::*:W:BW:"),
	(0,     0,     1,     'B',     2,     0, "WBW:::B::::W:BW:"),
	(0,     0,     1,     'B',     1,     0, "WBB:::B::::W:BW:"),
	(0,     1,     0,     'W',     9,     0, "WBB:::B::::W:BW:"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     0, ":::::::::::::W::"),
	(0,     0,     0,     '*',     7,     0, ":::::::::::::B::"),
	(0,     0,     1,     'W',     5,     0, ":::::::::::::B::"),
	(0,     0,     0,     ':',     14,     0, ":::::W:::::::B::"),
	(0,     0,     0,     ':',     6,     0, ":::::W:::::::B::"),
	(0,     0,     0,     'W',     7,     0, ":::::W:::::::B::"),
	(0,     0,     0,     ':',     7,     0, ":::::W:::::::B::"),
	(0,     0,     1,     '*',     9,     0, ":::::W:::::::B::"),
	(0,     0,     0,     'B',     11,     0, ":::::W:::*:::B::"),
	(0,     0,     1,     '*',     2,     0, ":::::W:::*:::B::"),
	(0,     0,     0,     '*',     13,     0, "::*::W:::*:::B::"),
	(0,     0,     0,     'W',     14,     0, "::*::W:::*:::B::"),
	(0,     0,     0,     '*',     9,     0, "::*::W:::*:::B::"),
	(0,     0,     0,     'B',     5,     0, "::*::W:::*:::B::"),
	(0,     0,     1,     'B',     14,     0, "::*::W:::*:::B::"),
	(0,     0,     0,     'B',     9,     0, "::*::W:::*:::BB:"),
	(0,     0,     1,     'B',     4,     0, "::*::W:::*:::BB:"),
	(0,     0,     1,     'W',     14,     0, "::*:BW:::*:::BB:"),
	(0,     0,     0,     '*',     7,     0, "::*:BW:::*:::BW:"),
	(0,     0,     1,     ':',     14,     0, "::*:BW:::*:::BW:"),
	(0,     0,     0,     ':',     5,     0, "::*:BW:::*:::BW:"),
	(0,     0,     0,     'W',     8,     0, "::*:BW:::*:::BW:"),
	(0,     0,     1,     ':',     14,     0, "::*:BW:::*:::BW:"),
	(0,     0,     0,     ':',     1,     0, "::*:BW:::*:::BW:"),
	(0,     1,     1,     'W',     6,     0, "::*:BW:::*:::BW:"),
	(0,     0,     1,     '*',     4,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     12,     0, "::::*:W:::::::::"),
	(0,     0,     0,     'B',     12,     0, "::::*:W:::::::::"),
	(0,     0,     0,     ':',     15,     0, "::::*:W:::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::*:W:::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::*:W:::::::::"),
	(0,     0,     1,     '*',     14,     0, "::*:*:W:::::::::"),
	(0,     1,     1,     '*',     2,     0, "::*:*:W:::::::*:"),
	(0,     0,     1,     'W',     5,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     6,     0, "::*::W::::::::::"),
	(0,     0,     1,     'W',     3,     0, "::*::W::::::::::"),
	(0,     0,     1,     'B',     15,     0, "::*W:W::::::::::"),
	(0,     1,     0,     'B',     13,     0, "::*W:W:::::::::B"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, "::::::::::W:::::"),
	(0,     0,     1,     'B',     2,     0, "::::::::::W:::::"),
	(0,     1,     0,     '*',     15,     0, "::B:::::::W:::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     10,     0, "::::::::::::::B:"),
	(0,     0,     0,     'W',     7,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     6,     0, "::::::::::::::B:"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::::B:"),
	(0,     0,     1,     'B',     13,     0, "::::::::::::::B:"),
	(0,     0,     1,     '*',     3,     0, ":::::::::::::BB:"),
	(0,     1,     0,     ':',     14,     0, ":::*:::::::::BB:"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     8,     0, "B::::W::::::::::"),
	(0,     0,     0,     'B',     7,     0, "B::::W::W:::::::"),
	(0,     0,     0,     'B',     15,     0, "B::::W::W:::::::"),
	(0,     0,     1,     'B',     4,     0, "B::::W::W:::::::"),
	(0,     0,     1,     'W',     9,     0, "B:::BW::W:::::::"),
	(0,     0,     0,     'B',     9,     0, "B:::BW::WW::::::"),
	(0,     0,     1,     '*',     14,     0, "B:::BW::WW::::::"),
	(0,     0,     0,     ':',     4,     0, "B:::BW::WW::::*:"),
	(0,     0,     1,     'B',     10,     0, "B:::BW::WW::::*:"),
	(0,     0,     0,     '*',     12,     0, "B:::BW::WWB:::*:"),
	(0,     1,     0,     '*',     10,     0, "B:::BW::WWB:::*:"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::::::W::::::::"),
	(0,     0,     1,     'W',     5,     0, ":::::::W::::::::"),
	(0,     0,     0,     'W',     13,     0, ":::::W:W::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::::W:W::::::::"),
	(0,     0,     1,     '*',     4,     0, ":::::W:W::::::W:"),
	(0,     0,     0,     '*',     0,     0, "::::*W:W::::::W:"),
	(0,     0,     1,     '*',     1,     0, "::::*W:W::::::W:"),
	(0,     0,     0,     'B',     11,     0, ":*::*W:W::::::W:"),
	(0,     0,     0,     ':',     2,     0, ":*::*W:W::::::W:"),
	(0,     0,     1,     'W',     5,     0, ":*::*W:W::::::W:"),
	(0,     0,     1,     'W',     4,     0, ":*::*W:W::::::W:"),
	(0,     0,     1,     ':',     15,     0, ":*::WW:W::::::W:"),
	(0,     0,     1,     ':',     0,     0, ":*::WW:W::::::W:"),
	(0,     0,     0,     'B',     7,     0, ":*::WW:W::::::W:"),
	(0,     0,     0,     'B',     11,     0, ":*::WW:W::::::W:"),
	(0,     0,     0,     '*',     7,     0, ":*::WW:W::::::W:"),
	(0,     0,     0,     '*',     15,     0, ":*::WW:W::::::W:"),
	(0,     0,     0,     ':',     0,     0, ":*::WW:W::::::W:"),
	(0,     0,     1,     ':',     4,     0, ":*::WW:W::::::W:"),
	(0,     0,     1,     ':',     8,     0, ":*::WW:W::::::W:"),
	(0,     0,     1,     'B',     0,     0, ":*::WW:W::::::W:"),
	(0,     0,     0,     ':',     15,     0, "B*::WW:W::::::W:"),
	(0,     0,     1,     'B',     0,     0, "B*::WW:W::::::W:"),
	(0,     0,     0,     ':',     2,     0, "B*::WW:W::::::W:"),
	(0,     0,     1,     '*',     12,     0, "B*::WW:W::::::W:"),
	(0,     1,     0,     '*',     0,     0, "B*::WW:W::::*:W:"),
	(0,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     0, ":::::::::::::*::"),
	(0,     0,     1,     'B',     14,     0, ":::::::::::::*::"),
	(0,     0,     0,     'W',     13,     0, ":::::::::::::*B:"),
	(0,     0,     1,     '*',     6,     0, ":::::::::::::*B:"),
	(0,     0,     0,     ':',     13,     0, "::::::*::::::*B:"),
	(0,     0,     0,     'B',     8,     0, "::::::*::::::*B:"),
	(0,     0,     0,     'B',     15,     0, "::::::*::::::*B:"),
	(0,     1,     0,     'B',     2,     0, "::::::*::::::*B:"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(1,     0,     0,     ':',     8,     0, ":::W::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     11,     0, "::::::::::::::B:"),
	(0,     0,     1,     'B',     0,     0, ":::::::::::B::::"),
	(0,     1,     0,     ':',     9,     0, "B::::::::::B::::"),
	(0,     1,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     11,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     4,     0, "::::::::::::W:::"),
	(0,     0,     1,     ':',     0,     0, "::::W:::::::W:::"),
	(0,     0,     1,     ':',     12,     0, "::::W:::::::W:::"),
	(0,     0,     1,     ':',     2,     0, "::::W:::::::W:::"),
	(0,     0,     0,     '*',     1,     0, "::::W:::::::W:::"),
	(0,     0,     0,     'W',     8,     0, "::::W:::::::W:::"),
	(0,     0,     1,     'W',     13,     0, "::::W:::::::W:::"),
	(0,     0,     0,     'B',     5,     0, "::::W:::::::WW::"),
	(0,     1,     1,     'B',     7,     0, "::::W:::::::WW::"),
	(0,     1,     1,     ':',     13,     0, ":::::::B::::::::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "::::::::*:::::::"),
	(0,     0,     1,     'W',     13,     0, "::::::::*:::*:::"),
	(0,     0,     1,     'W',     2,     0, "::::::::*:::*W::"),
	(0,     0,     1,     'W',     2,     0, "::W:::::*:::*W::"),
	(0,     0,     1,     ':',     2,     0, "::W:::::*:::*W::"),
	(0,     0,     1,     ':',     6,     0, "::W:::::*:::*W::"),
	(0,     0,     1,     'B',     8,     0, "::W:::::*:::*W::"),
	(0,     0,     1,     'W',     11,     0, "::W:::::B:::*W::"),
	(0,     0,     1,     '*',     8,     0, "::W:::::B::W*W::"),
	(0,     0,     0,     'W',     11,     0, "::W:::::W::W*W::"),
	(0,     0,     0,     'W',     15,     0, "::W:::::W::W*W::"),
	(0,     0,     1,     'B',     15,     0, "::W:::::W::W*W::"),
	(0,     0,     0,     'W',     6,     0, "::W:::::W::W*W:B"),
	(0,     0,     0,     '*',     4,     0, "::W:::::W::W*W:B"),
	(0,     0,     1,     'B',     8,     0, "::W:::::W::W*W:B"),
	(0,     0,     1,     'B',     0,     0, "::W:::::B::W*W:B"),
	(0,     0,     1,     'B',     0,     0, "B:W:::::B::W*W:B"),
	(0,     0,     1,     'W',     8,     0, "B:W:::::B::W*W:B"),
	(0,     1,     0,     '*',     2,     0, "B:W:::::W::W*W:B"),
	(1,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     6,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     4,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     15,     0, ":::::::::*::::::"),
	(0,     0,     0,     '*',     2,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     8,     0, ":::::::::*::::::"),
	(0,     0,     1,     'B',     5,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     4,     0, ":::::B:::*::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::B:::*::::::"),
	(0,     0,     0,     '*',     8,     0, ":::::B:::*::::::"),
	(0,     0,     0,     'B',     6,     0, ":::::B:::*::::::"),
	(0,     0,     1,     '*',     0,     0, ":::::B:::*::::::"),
	(0,     0,     1,     '*',     2,     0, "*::::B:::*::::::"),
	(0,     0,     0,     'W',     2,     0, "*:*::B:::*::::::"),
	(0,     0,     1,     '*',     10,     0, "*:*::B:::*::::::"),
	(0,     0,     1,     'W',     3,     0, "*:*::B:::**:::::"),
	(0,     0,     0,     'B',     3,     0, "*:*W:B:::**:::::"),
	(0,     0,     1,     ':',     7,     0, "*:*W:B:::**:::::"),
	(0,     0,     0,     'B',     14,     0, "*:*W:B:::**:::::"),
	(0,     1,     1,     ':',     10,     0, "*:*W:B:::**:::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     6,     0, "::::::W::::::::*"),
	(0,     0,     1,     '*',     5,     0, "::::::W::::::::*"),
	(0,     0,     0,     'W',     12,     0, ":::::*W::::::::*"),
	(0,     0,     1,     'B',     0,     0, ":::::*W::::::::*"),
	(0,     0,     0,     'W',     12,     0, "B::::*W::::::::*"),
	(0,     0,     0,     'W',     0,     0, "B::::*W::::::::*"),
	(0,     0,     1,     'B',     13,     0, "B::::*W::::::::*"),
	(0,     0,     0,     'B',     13,     0, "B::::*W::::::B:*"),
	(0,     0,     0,     'B',     11,     0, "B::::*W::::::B:*"),
	(0,     0,     1,     'B',     10,     0, "B::::*W::::::B:*"),
	(0,     0,     1,     ':',     11,     0, "B::::*W:::B::B:*"),
	(0,     0,     0,     '*',     7,     0, "B::::*W:::B::B:*"),
	(0,     0,     0,     'B',     9,     0, "B::::*W:::B::B:*"),
	(0,     0,     1,     '*',     8,     0, "B::::*W:::B::B:*"),
	(0,     0,     1,     'B',     6,     0, "B::::*W:*:B::B:*"),
	(0,     0,     0,     'B',     7,     0, "B::::*B:*:B::B:*"),
	(0,     0,     0,     ':',     0,     0, "B::::*B:*:B::B:*"),
	(0,     0,     0,     'B',     4,     0, "B::::*B:*:B::B:*"),
	(0,     0,     0,     '*',     1,     0, "B::::*B:*:B::B:*"),
	(0,     0,     0,     ':',     0,     0, "B::::*B:*:B::B:*"),
	(0,     0,     1,     'B',     9,     0, "B::::*B:*:B::B:*"),
	(0,     0,     0,     'W',     15,     0, "B::::*B:*BB::B:*"),
	(0,     0,     0,     '*',     6,     0, "B::::*B:*BB::B:*"),
	(0,     0,     1,     'B',     6,     0, "B::::*B:*BB::B:*"),
	(0,     0,     1,     ':',     14,     0, "B::::*B:*BB::B:*"),
	(0,     0,     1,     '*',     0,     0, "B::::*B:*BB::B:*"),
	(0,     1,     1,     'B',     7,     0, "W::::*B:*BB::B:*"),
	(0,     0,     1,     ':',     13,     0, ":::::::B::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::::B::::::::"),
	(0,     0,     1,     'W',     12,     0, ":::::::B::::::::"),
	(0,     0,     1,     'B',     3,     0, ":::::::B::::W:::"),
	(0,     0,     1,     'W',     12,     0, ":::B:::B::::W:::"),
	(0,     0,     0,     '*',     15,     0, ":::B:::B::::W:::"),
	(0,     0,     1,     'W',     1,     0, ":::B:::B::::W:::"),
	(0,     0,     0,     '*',     5,     0, ":W:B:::B::::W:::"),
	(0,     0,     1,     'W',     7,     0, ":W:B:::B::::W:::"),
	(0,     0,     1,     ':',     11,     0, ":W:B:::W::::W:::"),
	(0,     0,     0,     'B',     8,     0, ":W:B:::W::::W:::"),
	(0,     0,     1,     'B',     1,     0, ":W:B:::W::::W:::"),
	(0,     0,     0,     'W',     14,     0, ":B:B:::W::::W:::"),
	(0,     0,     0,     '*',     4,     0, ":B:B:::W::::W:::"),
	(0,     1,     1,     ':',     5,     0, ":B:B:::W::::W:::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     0, ":::W::::::::::::"),
	(0,     0,     0,     'W',     8,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     11,     0, ":::W::::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::W::::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::W::::::::::::"),
	(0,     1,     0,     'W',     3,     0, ":::W::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     11,     0, ":::::W::::*:::::"),
	(0,     0,     0,     '*',     4,     0, ":::::W::::*:::::"),
	(0,     0,     1,     ':',     0,     0, ":::::W::::*:::::"),
	(0,     0,     0,     '*',     12,     0, ":::::W::::*:::::"),
	(0,     0,     1,     'B',     3,     0, ":::::W::::*:::::"),
	(0,     0,     1,     'B',     15,     0, ":::B:W::::*:::::"),
	(0,     0,     0,     'B',     15,     0, ":::B:W::::*::::B"),
	(0,     0,     1,     'B',     7,     0, ":::B:W::::*::::B"),
	(0,     0,     1,     ':',     9,     0, ":::B:W:B::*::::B"),
	(0,     0,     0,     ':',     7,     0, ":::B:W:B::*::::B"),
	(0,     1,     0,     'W',     0,     0, ":::B:W:B::*::::B"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     13,     0, ":*:::::::::B::::"),
	(0,     1,     1,     ':',     5,     0, ":*:::::::::B::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, ":::::::::::B::::"),
	(0,     1,     1,     ':',     8,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     8,     0, ":::B::::::::::::"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     7,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, "::W:::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::W:::::::::::::"),
	(0,     0,     0,     'B',     1,     0, "::W:::::::::::::"),
	(0,     0,     0,     'B',     11,     0, "::W:::::::::::::"),
	(0,     0,     0,     'B',     14,     0, "::W:::::::::::::"),
	(0,     0,     1,     'W',     3,     0, "::W:::::::::::::"),
	(0,     0,     0,     ':',     1,     0, "::WW::::::::::::"),
	(0,     0,     1,     '*',     7,     0, "::WW::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::WW:::*::::::::"),
	(0,     0,     0,     'B',     7,     0, "::WW:::*::::::::"),
	(0,     0,     0,     ':',     13,     0, "::WW:::*::::::::"),
	(0,     0,     1,     'B',     9,     0, "::WW:::*::::::::"),
	(0,     0,     0,     'W',     10,     0, "::WW:::*:B::::::"),
	(0,     0,     1,     'B',     4,     0, "::WW:::*:B::::::"),
	(0,     0,     0,     'W',     14,     0, "::WWB::*:B::::::"),
	(0,     0,     0,     ':',     6,     0, "::WWB::*:B::::::"),
	(0,     0,     1,     'W',     11,     0, "::WWB::*:B::::::"),
	(0,     0,     1,     '*',     1,     0, "::WWB::*:B:W::::"),
	(0,     0,     0,     '*',     7,     0, ":*WWB::*:B:W::::"),
	(0,     0,     1,     ':',     9,     0, ":*WWB::*:B:W::::"),
	(0,     0,     1,     'W',     4,     0, ":*WWB::*:B:W::::"),
	(0,     1,     1,     'B',     11,     0, ":*WWW::*:B:W::::"),
	(0,     0,     1,     '*',     13,     0, ":::::::::::B::::"),
	(0,     0,     1,     ':',     10,     0, ":::::::::::B:*::"),
	(0,     0,     0,     '*',     10,     0, ":::::::::::B:*::"),
	(0,     0,     1,     ':',     15,     0, ":::::::::::B:*::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::B:*::"),
	(0,     0,     0,     'W',     11,     0, ":::::::::::B:*::"),
	(0,     0,     0,     '*',     4,     0, ":::::::::::B:*::"),
	(1,     0,     0,     'B',     1,     0, ":::::::::::B:*::"),
	(0,     1,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, ":::::::::::::::*"),
	(0,     1,     0,     'W',     7,     0, ":::::::::::::::*"),
	(0,     0,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     0, "::::B:::::::::::"),
	(0,     0,     0,     'B',     10,     0, "::::B:::::::::*:"),
	(0,     0,     1,     '*',     14,     0, "::::B:::::::::*:"),
	(0,     0,     0,     'W',     13,     0, "::::B:::::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::B:::::::::::"),
	(0,     0,     1,     'W',     12,     0, "::::B:::::::::::"),
	(0,     0,     0,     ':',     2,     0, "::::B:::::::W:::"),
	(0,     0,     0,     '*',     4,     0, "::::B:::::::W:::"),
	(0,     0,     0,     'B',     4,     0, "::::B:::::::W:::"),
	(0,     0,     0,     ':',     15,     0, "::::B:::::::W:::"),
	(0,     0,     0,     'W',     11,     0, "::::B:::::::W:::"),
	(0,     0,     0,     ':',     1,     0, "::::B:::::::W:::"),
	(0,     1,     0,     ':',     4,     0, "::::B:::::::W:::"),
	(0,     1,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     0,     1, "::::::::::::::::"),
	(1,     0,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     0, "::B:::::::::::::"),
	(0,     0,     1,     ':',     8,     0, "::B:*:::::::::::"),
	(0,     0,     0,     'B',     9,     0, "::B:*:::::::::::"),
	(0,     0,     1,     'W',     12,     0, "::B:*:::::::::::"),
	(0,     0,     0,     'B',     5,     0, "::B:*:::::::W:::"),
	(0,     0,     0,     'B',     6,     0, "::B:*:::::::W:::"),
	(0,     0,     0,     '*',     9,     0, "::B:*:::::::W:::"),
	(0,     0,     0,     '*',     5,     0, "::B:*:::::::W:::"),
	(0,     0,     1,     '*',     2,     0, "::B:*:::::::W:::"),
	(0,     0,     1,     ':',     12,     0, "::W:*:::::::W:::"),
	(0,     0,     1,     '*',     4,     0, "::W:*:::::::W:::"),
	(0,     0,     0,     'B',     1,     0, "::W:::::::::W:::"),
	(0,     1,     0,     '*',     13,     0, "::W:::::::::W:::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, "::::W:::::::::::"),
	(0,     0,     0,     'B',     9,     0, "::::W:::::::::::"),
	(0,     1,     0,     'B',     12,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     0, "B:::::::::::::::"),
	(0,     0,     0,     'W',     3,     0, "B:B:::::::::::::"),
	(0,     0,     0,     'B',     3,     0, "B:B:::::::::::::"),
	(0,     0,     1,     'W',     13,     0, "B:B:::::::::::::"),
	(1,     0,     1,     'W',     7,     0, "B:B::::::::::W::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     0, "::::B:::::::::::"),
	(1,     0,     0,     '*',     9,     0, "::::B::::*::::::"),
	(0,     0,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     0, "::::::::W:::::::"),
	(0,     0,     0,     'W',     3,     0, "::::*:::W:::::::"),
	(0,     0,     1,     'W',     13,     0, "::::*:::W:::::::"),
	(0,     0,     1,     '*',     4,     0, "::::*:::W::::W::"),
	(0,     1,     0,     '*',     7,     0, "::::::::W::::W::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     0, "::::::::B:::::::"),
	(0,     0,     0,     '*',     1,     0, "::::::::B:::::::"),
	(0,     0,     0,     'B',     14,     0, "::::::::B:::::::"),
	(0,     1,     1,     'W',     5,     0, "::::::::B:::::::"),
	(0,     0,     0,     'B',     12,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     11,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     0,     0, ":::::W::::::::::"),
	(0,     1,     0,     ':',     13,     0, "W::::W::::::::::"),
	(1,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     0, ":::W::::::::::::"),
	(0,     0,     1,     'B',     1,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     3,     0, ":B:W::::::::::::"),
	(1,     0,     0,     '*',     6,     0, ":B:W::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     14,     0, "B:::::::::::::::"),
	(0,     1,     0,     ':',     15,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     4,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::::::B::::::::"),
	(0,     0,     1,     'B',     13,     0, ":::::::B::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::::::B:::::B::"),
	(0,     0,     0,     '*',     7,     0, ":::::::B:::::B::"),
	(0,     0,     1,     'B',     13,     0, ":::::::B:::::B::"),
	(0,     0,     0,     '*',     5,     0, ":::::::B:::::B::"),
	(0,     0,     0,     ':',     0,     0, ":::::::B:::::B::"),
	(0,     0,     0,     ':',     1,     0, ":::::::B:::::B::"),
	(0,     0,     0,     'W',     7,     0, ":::::::B:::::B::"),
	(0,     0,     0,     '*',     3,     0, ":::::::B:::::B::"),
	(0,     0,     1,     '*',     6,     0, ":::::::B:::::B::"),
	(0,     0,     1,     ':',     15,     0, "::::::*B:::::B::"),
	(0,     0,     0,     ':',     9,     0, "::::::*B:::::B::"),
	(0,     0,     1,     'W',     9,     0, "::::::*B:::::B::"),
	(0,     0,     1,     'W',     2,     0, "::::::*B:W:::B::"),
	(0,     1,     0,     'B',     3,     0, "::W:::*B:W:::B::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     0, ":W::::::::::::::"),
	(0,     0,     1,     '*',     4,     0, ":W::::::::::::*:"),
	(0,     1,     1,     'W',     4,     0, ":W::*:::::::::*:"),
	(0,     0,     1,     '*',     13,     0, "::::W:::::::::::"),
	(0,     0,     1,     ':',     4,     0, "::::W::::::::*::"),
	(0,     0,     1,     '*',     1,     0, "::::W::::::::*::"),
	(0,     0,     1,     'B',     3,     0, ":*::W::::::::*::"),
	(0,     0,     1,     '*',     15,     0, ":*:BW::::::::*::"),
	(0,     0,     0,     '*',     12,     0, ":*:BW::::::::*:*"),
	(0,     0,     0,     ':',     0,     0, ":*:BW::::::::*:*"),
	(0,     0,     0,     'B',     9,     0, ":*:BW::::::::*:*"),
	(0,     0,     1,     ':',     9,     0, ":*:BW::::::::*:*"),
	(0,     0,     1,     ':',     1,     0, ":*:BW::::::::*:*"),
	(0,     0,     0,     'W',     8,     0, ":*:BW::::::::*:*"),
	(0,     0,     1,     'W',     6,     0, ":*:BW::::::::*:*"),
	(1,     0,     1,     '*',     9,     0, ":*:BW:W::::::*:*"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     3,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     15,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     1,     0, "::::::*::::::::*"),
	(0,     0,     0,     '*',     11,     0, ":*::::*::::::::*"),
	(0,     1,     0,     '*',     12,     0, ":*::::*::::::::*"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     6,     0, ":B::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     0, "B:::::::::::::::"),
	(1,     0,     1,     'W',     5,     0, "B::::::::::::B::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     0, "::*:::::::::::::"),
	(0,     0,     1,     '*',     4,     0, "::*:::::::::::::"),
	(0,     1,     0,     ':',     2,     0, "::*:*:::::::::::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::::::B:::::::"),
	(0,     0,     1,     'W',     6,     0, "::*:::::B:::::::"),
	(0,     0,     1,     '*',     13,     0, "::*:::W:B:::::::"),
	(0,     0,     1,     ':',     14,     0, "::*:::W:B::::*::"),
	(0,     0,     1,     'W',     11,     0, "::*:::W:B::::*::"),
	(0,     0,     0,     ':',     14,     0, "::*:::W:B::W:*::"),
	(0,     0,     0,     'B',     9,     0, "::*:::W:B::W:*::"),
	(0,     0,     1,     'B',     13,     0, "::*:::W:B::W:*::"),
	(0,     0,     0,     'B',     11,     0, "::*:::W:B::W:B::"),
	(0,     0,     1,     'B',     6,     0, "::*:::W:B::W:B::"),
	(0,     0,     0,     ':',     3,     0, "::*:::B:B::W:B::"),
	(0,     0,     1,     'W',     10,     0, "::*:::B:B::W:B::"),
	(0,     0,     0,     'W',     7,     0, "::*:::B:B:WW:B::"),
	(0,     0,     0,     ':',     3,     0, "::*:::B:B:WW:B::"),
	(0,     0,     1,     'W',     3,     0, "::*:::B:B:WW:B::"),
	(0,     0,     1,     '*',     3,     0, "::*W::B:B:WW:B::"),
	(0,     0,     1,     '*',     0,     0, "::*B::B:B:WW:B::"),
	(0,     0,     0,     '*',     2,     0, "*:*B::B:B:WW:B::"),
	(0,     1,     1,     'B',     12,     0, "*:*B::B:B:WW:B::"),
	(0,     0,     1,     ':',     15,     0, "::::::::::::B:::"),
	(0,     0,     0,     ':',     14,     0, "::::::::::::B:::"),
	(0,     1,     1,     'B',     15,     0, "::::::::::::B:::"),
	(0,     0,     0,     '*',     8,     0, ":::::::::::::::B"),
	(0,     0,     1,     '*',     11,     0, ":::::::::::::::B"),
	(0,     0,     0,     ':',     15,     0, ":::::::::::*:::B"),
	(0,     0,     0,     ':',     7,     0, ":::::::::::*:::B"),
	(0,     0,     0,     'B',     2,     0, ":::::::::::*:::B"),
	(0,     0,     0,     'W',     9,     0, ":::::::::::*:::B"),
	(0,     0,     0,     '*',     7,     0, ":::::::::::*:::B"),
	(0,     1,     1,     '*',     8,     0, ":::::::::::*:::B"),
	(0,     0,     1,     ':',     11,     0, "::::::::*:::::::"),
	(0,     0,     0,     'W',     9,     0, "::::::::*:::::::"),
	(0,     0,     0,     'W',     15,     0, "::::::::*:::::::"),
	(0,     0,     1,     '*',     8,     0, "::::::::*:::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     9,     0, "::::::*:::::::::"),
	(0,     0,     0,     ':',     2,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     1,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     12,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     15,     0, "::::::*:::::*:::"),
	(0,     0,     1,     ':',     11,     0, "::::::*:::::*:::"),
	(0,     0,     1,     ':',     5,     0, "::::::*:::::*:::"),
	(0,     0,     0,     '*',     13,     0, "::::::*:::::*:::"),
	(0,     1,     1,     ':',     11,     0, "::::::*:::::*:::"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     9,     0, "::::::B::::::::B"),
	(0,     1,     1,     '*',     14,     0, "::::::B::::::::B"),
	(0,     1,     0,     ':',     3,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     3,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::::::*"),
	(0,     0,     1,     'B',     2,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     7,     0, "::B::::::::::::*"),
	(0,     0,     0,     'W',     9,     0, "::B::::::::::::*"),
	(0,     0,     1,     '*',     3,     0, "::B::::::::::::*"),
	(0,     0,     1,     ':',     8,     0, "::B*:::::::::::*"),
	(0,     0,     0,     '*',     13,     0, "::B*:::::::::::*"),
	(0,     0,     0,     'B',     1,     0, "::B*:::::::::::*"),
	(0,     0,     0,     '*',     4,     0, "::B*:::::::::::*"),
	(0,     0,     1,     '*',     15,     0, "::B*:::::::::::*"),
	(0,     0,     1,     '*',     5,     0, "::B*::::::::::::"),
	(0,     0,     0,     'B',     13,     0, "::B*:*::::::::::"),
	(0,     1,     1,     'B',     8,     0, "::B*:*::::::::::"),
	(0,     1,     0,     'B',     3,     0, "::::::::B:::::::"),
	(1,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     6,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::::*:::::::::"),
	(0,     0,     0,     'W',     11,     0, "::*:::*:::::::::"),
	(0,     0,     0,     '*',     0,     0, "::*:::*:::::::::"),
	(0,     0,     0,     'B',     14,     0, "::*:::*:::::::::"),
	(0,     0,     1,     '*',     11,     0, "::*:::*:::::::::"),
	(0,     1,     0,     'B',     11,     0, "::*:::*::::*::::"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::*::::::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     6,     0, ":::*::::::::::::"),
	(0,     0,     1,     '*',     2,     0, ":::*::::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::**::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "::**::::::::::::"),
	(0,     0,     1,     'B',     13,     0, "::**::::::::*:::"),
	(0,     0,     1,     ':',     15,     0, "::**::::::::*B::"),
	(0,     0,     0,     'W',     5,     0, "::**::::::::*B::"),
	(0,     0,     1,     ':',     3,     0, "::**::::::::*B::"),
	(0,     0,     1,     'B',     5,     0, "::**::::::::*B::"),
	(0,     0,     1,     'W',     14,     0, "::**:B::::::*B::"),
	(0,     0,     1,     '*',     1,     0, "::**:B::::::*BW:"),
	(0,     0,     0,     '*',     2,     0, ":***:B::::::*BW:"),
	(1,     0,     1,     '*',     6,     0, ":***:B::::::*BW:"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     0, ":B::::::::::::::"),
	(0,     1,     0,     '*',     1,     0, ":B::::*:::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     0,     0, "::::::W::W::::::"),
	(0,     0,     1,     ':',     10,     0, "::::::W::W::::::"),
	(0,     0,     1,     '*',     5,     0, "::::::W::W::::::"),
	(0,     0,     1,     'W',     9,     0, ":::::*W::W::::::"),
	(0,     0,     1,     'B',     2,     0, ":::::*W::W::::::"),
	(0,     0,     1,     'B',     3,     0, "::B::*W::W::::::"),
	(0,     1,     0,     'W',     13,     0, "::BB:*W::W::::::"),
	(0,     1,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "W:::::::::::::::"),
	(0,     0,     0,     '*',     7,     0, "W:::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, "W:::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, "W::::::::::B::::"),
	(0,     0,     0,     ':',     13,     0, "W::::::::::W::::"),
	(0,     0,     0,     ':',     4,     0, "W::::::::::W::::"),
	(0,     0,     0,     '*',     7,     0, "W::::::::::W::::"),
	(0,     0,     0,     'B',     15,     0, "W::::::::::W::::"),
	(0,     1,     0,     'B',     10,     0, "W::::::::::W::::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     12,     0, ":::::::*::::::::"),
	(0,     0,     1,     'B',     2,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     5,     0, "::B:::::::::W:::"),
	(0,     0,     1,     'B',     7,     0, "::B:::::::::W:::"),
	(0,     0,     1,     '*',     0,     0, "::B::::B::::W:::"),
	(0,     0,     0,     'B',     15,     0, "*:B::::B::::W:::"),
	(0,     0,     0,     'W',     4,     0, "*:B::::B::::W:::"),
	(0,     0,     1,     'B',     15,     0, "*:B::::B::::W:::"),
	(0,     0,     0,     ':',     5,     0, "*:B::::B::::W::B"),
	(0,     0,     0,     '*',     7,     0, "*:B::::B::::W::B"),
	(0,     0,     0,     ':',     12,     0, "*:B::::B::::W::B"),
	(0,     1,     1,     'W',     8,     0, "*:B::::B::::W::B"),
	(0,     0,     0,     '*',     11,     0, "::::::::W:::::::"),
	(0,     0,     1,     ':',     7,     0, "::::::::W:::::::"),
	(0,     0,     1,     ':',     6,     0, "::::::::W:::::::"),
	(0,     0,     1,     'W',     11,     0, "::::::::W:::::::"),
	(0,     0,     1,     '*',     0,     0, "::::::::W::W::::"),
	(0,     0,     1,     'B',     8,     0, "*:::::::W::W::::"),
	(0,     0,     1,     '*',     14,     0, "*:::::::B::W::::"),
	(0,     0,     0,     '*',     15,     0, "*:::::::B::W::*:"),
	(0,     0,     0,     ':',     11,     0, "*:::::::B::W::*:"),
	(0,     0,     0,     'W',     1,     0, "*:::::::B::W::*:"),
	(0,     1,     1,     '*',     5,     0, "*:::::::B::W::*:"),
	(0,     0,     1,     'B',     10,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::::*::::B:::::"),
	(0,     0,     1,     '*',     5,     0, ":::::*::::B:::::"),
	(0,     0,     1,     ':',     15,     0, "::::::::::B:::::"),
	(0,     0,     1,     'B',     7,     0, "::::::::::B:::::"),
	(0,     0,     1,     '*',     7,     0, ":::::::B::B:::::"),
	(0,     0,     1,     ':',     9,     0, ":::::::W::B:::::"),
	(0,     1,     0,     ':',     11,     0, ":::::::W::B:::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     11,     0, ":::::::::*::::::"),
	(0,     0,     0,     '*',     3,     0, ":::::::::*:*::::"),
	(0,     0,     1,     'B',     15,     0, ":::::::::*:*::::"),
	(0,     1,     1,     'B',     5,     0, ":::::::::*:*:::B"),
	(0,     0,     1,     '*',     5,     0, ":::::B::::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     5,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::WW:::::::::"),
	(0,     0,     0,     'B',     3,     0, ":::::WW:::::::::"),
	(0,     1,     0,     ':',     2,     0, ":::::WW:::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, ":::::W::::::::::"),
	(0,     0,     1,     '*',     15,     0, ":::::W:::W::::::"),
	(0,     0,     0,     ':',     0,     0, ":::::W:::W:::::*"),
	(0,     1,     1,     '*',     2,     0, ":::::W:::W:::::*"),
	(0,     0,     0,     'B',     7,     0, "::*:::::::::::::"),
	(0,     0,     1,     '*',     10,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     10,     0, "::*:::::::*:::::"),
	(0,     0,     0,     'W',     0,     0, "::*:::::::B:::::"),
	(0,     0,     0,     'B',     1,     0, "::*:::::::B:::::"),
	(0,     0,     0,     'W',     13,     0, "::*:::::::B:::::"),
	(0,     0,     0,     'B',     9,     0, "::*:::::::B:::::"),
	(1,     0,     0,     ':',     14,     0, "::*:::::::B:::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     0, ":::::B::::::::::"),
	(0,     0,     1,     'W',     5,     0, ":::::B::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::W::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":::::W::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":::::W::::::*:::"),
	(0,     1,     1,     ':',     14,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     12,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     0,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     7,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     15,     0, "::::::::::::::*:"),
	(0,     0,     1,     ':',     1,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     3,     0, "::::::::::::::*:"),
	(0,     0,     0,     ':',     2,     0, "::::::::::::::*:"),
	(0,     1,     0,     '*',     11,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     0, ":::*::::::::::::"),
	(0,     1,     0,     ':',     9,     0, ":::*::B:::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     2,     0, ":::::W::::::::::"),
	(0,     0,     1,     '*',     9,     0, "::W::W::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::W::W:::*::::::"),
	(0,     0,     0,     ':',     10,     0, "::W::W:::*::::::"),
	(0,     0,     0,     'B',     7,     0, "::W::W:::*::::::"),
	(0,     0,     0,     'B',     13,     0, "::W::W:::*::::::"),
	(0,     0,     1,     '*',     14,     0, "::W::W:::*::::::"),
	(0,     0,     0,     'W',     4,     0, "::W::W:::*::::*:"),
	(0,     0,     1,     ':',     13,     0, "::W::W:::*::::*:"),
	(0,     1,     0,     '*',     0,     0, "::W::W:::*::::*:"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     0, "::::::::::::B:::"),
	(0,     0,     1,     ':',     15,     0, "::::::::::::BW::"),
	(0,     0,     0,     'B',     13,     0, "::::::::::::BW::"),
	(0,     0,     0,     ':',     12,     0, "::::::::::::BW::"),
	(0,     0,     0,     'W',     9,     0, "::::::::::::BW::"),
	(0,     0,     0,     'B',     7,     0, "::::::::::::BW::"),
	(0,     1,     0,     'B',     5,     0, "::::::::::::BW::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     0, ":::*::::::::::::"),
	(0,     0,     1,     'W',     7,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":::*:::W::::::::"),
	(0,     0,     1,     ':',     9,     0, ":::*:::W::::::::"),
	(0,     0,     1,     '*',     0,     0, ":::*:::W::::::::"),
	(0,     0,     1,     ':',     1,     0, "*::*:::W::::::::"),
	(0,     0,     1,     '*',     11,     0, "*::*:::W::::::::"),
	(0,     0,     0,     ':',     7,     0, "*::*:::W:::*::::"),
	(0,     0,     0,     'W',     2,     0, "*::*:::W:::*::::"),
	(0,     0,     0,     'B',     15,     0, "*::*:::W:::*::::"),
	(0,     1,     0,     ':',     5,     0, "*::*:::W:::*::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     0, "::::::::::*:::::"),
	(0,     0,     1,     'W',     10,     0, "::::::::::*:::::"),
	(0,     1,     0,     'W',     1,     0, "::::::::::W:::::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::W::::::::::::"),
	(1,     0,     1,     ':',     13,     0, ":::W::::::::::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     2,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     10,     0, "::B::::::::B::::"),
	(0,     0,     0,     'W',     1,     0, "::B:::::::*B::::"),
	(0,     0,     0,     ':',     5,     0, "::B:::::::*B::::"),
	(0,     0,     1,     ':',     5,     0, "::B:::::::*B::::"),
	(0,     0,     1,     'B',     4,     0, "::B:::::::*B::::"),
	(0,     0,     1,     'B',     0,     0, "::B:B:::::*B::::"),
	(0,     0,     1,     ':',     12,     0, "B:B:B:::::*B::::"),
	(0,     0,     1,     'B',     15,     0, "B:B:B:::::*B::::"),
	(0,     0,     0,     ':',     5,     0, "B:B:B:::::*B:::B"),
	(0,     1,     1,     'W',     14,     0, "B:B:B:::::*B:::B"),
	(0,     1,     1,     'W',     7,     0, "::::::::::::::W:"),
	(0,     0,     1,     'B',     8,     0, ":::::::W::::::::"),
	(0,     0,     1,     'W',     4,     0, ":::::::WB:::::::"),
	(0,     0,     0,     'W',     6,     0, "::::W::WB:::::::"),
	(0,     0,     0,     'W',     11,     0, "::::W::WB:::::::"),
	(0,     1,     1,     'W',     4,     0, "::::W::WB:::::::"),
	(0,     0,     0,     'W',     5,     0, "::::W:::::::::::"),
	(0,     0,     0,     ':',     14,     0, "::::W:::::::::::"),
	(0,     0,     0,     'W',     13,     0, "::::W:::::::::::"),
	(0,     0,     1,     ':',     12,     0, "::::W:::::::::::"),
	(0,     0,     0,     ':',     13,     0, "::::W:::::::::::"),
	(0,     0,     0,     'W',     11,     0, "::::W:::::::::::"),
	(0,     0,     1,     ':',     0,     0, "::::W:::::::::::"),
	(0,     1,     1,     '*',     7,     0, "::::W:::::::::::"),
	(0,     0,     1,     'W',     9,     0, ":::::::*::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::::*:W::::::"),
	(0,     0,     1,     'B',     6,     0, ":::::::*:W::::::"),
	(0,     0,     0,     'W',     2,     0, "::::::B*:W::::::"),
	(0,     0,     1,     'B',     2,     0, "::::::B*:W::::::"),
	(0,     0,     1,     'W',     10,     0, "::B:::B*:W::::::"),
	(0,     1,     0,     'B',     2,     0, "::B:::B*:WW:::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     0,     0, "*:::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     1,     0, "*::::::::::::::W"),
	(0,     0,     1,     'B',     10,     0, "*::::::::::::::W"),
	(0,     0,     0,     ':',     1,     0, "*:::::::::B::::W"),
	(0,     0,     0,     '*',     13,     0, "*:::::::::B::::W"),
	(0,     0,     1,     'B',     8,     0, "*:::::::::B::::W"),
	(0,     0,     0,     'W',     4,     0, "*:::::::B:B::::W"),
	(0,     0,     0,     'B',     11,     0, "*:::::::B:B::::W"),
	(0,     0,     0,     'B',     14,     0, "*:::::::B:B::::W"),
	(0,     0,     0,     'B',     8,     0, "*:::::::B:B::::W"),
	(0,     0,     1,     '*',     1,     0, "*:::::::B:B::::W"),
	(0,     0,     1,     ':',     2,     0, "**::::::B:B::::W"),
	(0,     0,     0,     'B',     13,     0, "**::::::B:B::::W"),
	(0,     0,     0,     ':',     10,     0, "**::::::B:B::::W"),
	(0,     0,     0,     ':',     4,     0, "**::::::B:B::::W"),
	(0,     0,     0,     'W',     12,     0, "**::::::B:B::::W"),
	(0,     0,     1,     'B',     14,     0, "**::::::B:B::::W"),
	(0,     0,     1,     'B',     1,     0, "**::::::B:B:::BW"),
	(0,     0,     1,     '*',     8,     0, "*B::::::B:B:::BW"),
	(0,     0,     1,     'W',     10,     0, "*B::::::W:B:::BW"),
	(0,     0,     0,     ':',     1,     0, "*B::::::W:W:::BW"),
	(0,     0,     1,     'W',     9,     0, "*B::::::W:W:::BW"),
	(0,     0,     1,     'B',     4,     0, "*B::::::WWW:::BW"),
	(0,     0,     1,     'B',     5,     0, "*B::B:::WWW:::BW"),
	(0,     0,     0,     'W',     5,     0, "*B::BB::WWW:::BW"),
	(0,     0,     1,     'W',     1,     0, "*B::BB::WWW:::BW"),
	(0,     0,     1,     ':',     14,     0, "*W::BB::WWW:::BW"),
	(0,     0,     1,     'B',     6,     0, "*W::BB::WWW:::BW"),
	(0,     0,     0,     '*',     10,     0, "*W::BBB:WWW:::BW"),
	(0,     0,     0,     'B',     12,     0, "*W::BBB:WWW:::BW"),
	(0,     0,     0,     ':',     12,     0, "*W::BBB:WWW:::BW"),
	(0,     0,     1,     'W',     14,     0, "*W::BBB:WWW:::BW"),
	(0,     0,     1,     'B',     0,     0, "*W::BBB:WWW:::WW"),
	(0,     0,     0,     ':',     13,     0, "BW::BBB:WWW:::WW"),
	(0,     0,     1,     '*',     15,     0, "BW::BBB:WWW:::WW"),
	(0,     0,     1,     'B',     1,     0, "BW::BBB:WWW:::WB"),
	(0,     0,     0,     ':',     4,     0, "BB::BBB:WWW:::WB"),
	(0,     0,     1,     '*',     4,     0, "BB::BBB:WWW:::WB"),
	(0,     0,     1,     'B',     1,     0, "BB::WBB:WWW:::WB"),
	(0,     0,     0,     ':',     6,     0, "BB::WBB:WWW:::WB"),
	(0,     0,     1,     'B',     6,     0, "BB::WBB:WWW:::WB"),
	(0,     0,     0,     'W',     1,     0, "BB::WBB:WWW:::WB"),
	(0,     0,     0,     ':',     15,     0, "BB::WBB:WWW:::WB"),
	(0,     1,     0,     'B',     2,     0, "BB::WBB:WWW:::WB"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     6,     0, "::::::W:::::::W:"),
	(0,     0,     1,     'B',     2,     0, "::::::B:::::::W:"),
	(0,     0,     1,     'B',     15,     0, "::B:::B:::::::W:"),
	(0,     0,     0,     '*',     2,     0, "::B:::B:::::::WB"),
	(0,     0,     0,     ':',     8,     0, "::B:::B:::::::WB"),
	(0,     1,     1,     '*',     11,     0, "::B:::B:::::::WB"),
	(0,     0,     1,     '*',     8,     0, ":::::::::::*::::"),
	(0,     0,     0,     '*',     0,     0, "::::::::*::*::::"),
	(0,     1,     0,     'W',     15,     0, "::::::::*::*::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     0, "::::::::::::*:::"),
	(0,     0,     0,     'W',     6,     0, "::::::::::W:*:::"),
	(0,     0,     1,     'B',     4,     0, "::::::::::W:*:::"),
	(0,     0,     1,     '*',     6,     0, "::::B:::::W:*:::"),
	(0,     0,     1,     'B',     14,     0, "::::B:*:::W:*:::"),
	(0,     0,     1,     'W',     9,     0, "::::B:*:::W:*:B:"),
	(0,     0,     0,     '*',     4,     0, "::::B:*::WW:*:B:"),
	(0,     1,     0,     'W',     7,     0, "::::B:*::WW:*:B:"),
	(0,     0,     0,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     0, ":::B::::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":::B:::*::::::::"),
	(0,     0,     1,     'W',     0,     0, ":::B:::*::::::::"),
	(0,     1,     1,     'W',     6,     0, "W::B:::*::::::::"),
	(0,     0,     0,     '*',     2,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     3,     0, "::::::W:::::::::"),
	(0,     0,     0,     '*',     5,     0, "::::::W:::::::::"),
	(0,     1,     0,     'W',     4,     0, "::::::W:::::::::"),
	(1,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(1,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     6,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     11,     0, "::::::W:::::::B:"),
	(0,     0,     1,     '*',     6,     0, "::::::W::::W::B:"),
	(0,     0,     0,     ':',     12,     0, "::::::B::::W::B:"),
	(0,     0,     0,     'B',     11,     0, "::::::B::::W::B:"),
	(0,     0,     0,     '*',     15,     0, "::::::B::::W::B:"),
	(0,     1,     1,     ':',     11,     0, "::::::B::::W::B:"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, ":*::::::::::::::"),
	(0,     1,     0,     'W',     7,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     14,     0, "::::::::W:::::::"),
	(0,     1,     1,     'B',     12,     0, "::::::::::::::B:"),
	(0,     0,     1,     '*',     2,     0, "::::::::::::B:::"),
	(0,     0,     1,     'B',     14,     0, "::*:::::::::B:::"),
	(0,     0,     1,     ':',     1,     0, "::*:::::::::B:B:"),
	(0,     0,     1,     'B',     3,     0, "::*:::::::::B:B:"),
	(0,     0,     1,     'W',     11,     0, "::*B::::::::B:B:"),
	(0,     0,     1,     'W',     9,     0, "::*B:::::::WB:B:"),
	(0,     1,     1,     'B',     14,     0, "::*B:::::W:WB:B:"),
	(0,     0,     0,     'B',     4,     0, "::::::::::::::B:"),
	(0,     0,     0,     'W',     5,     0, "::::::::::::::B:"),
	(0,     0,     1,     'B',     11,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     6,     0, ":::::::::::B::B:"),
	(0,     0,     0,     'W',     8,     0, ":::::::::::B::B:"),
	(0,     0,     1,     '*',     6,     0, ":::::::::::B::B:"),
	(0,     0,     0,     'W',     0,     0, "::::::*::::B::B:"),
	(0,     0,     0,     'B',     11,     0, "::::::*::::B::B:"),
	(0,     0,     0,     '*',     0,     0, "::::::*::::B::B:"),
	(0,     0,     1,     ':',     0,     0, "::::::*::::B::B:"),
	(0,     0,     1,     ':',     10,     0, "::::::*::::B::B:"),
	(0,     1,     1,     'B',     3,     0, "::::::*::::B::B:"),
	(0,     0,     0,     '*',     7,     0, ":::B::::::::::::"),
	(0,     0,     0,     '*',     6,     0, ":::B::::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":::B::::::::::::"),
	(0,     0,     0,     'B',     4,     0, ":::B::W:::::::::"),
	(0,     0,     0,     '*',     2,     0, ":::B::W:::::::::"),
	(0,     0,     0,     'W',     14,     0, ":::B::W:::::::::"),
	(0,     0,     1,     'B',     9,     0, ":::B::W:::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::B::W::B::::::"),
	(0,     0,     0,     'W',     8,     0, ":::B::W::B::::::"),
	(0,     0,     1,     'W',     7,     0, ":::B::W::B::::::"),
	(0,     0,     1,     ':',     1,     0, ":::B::WW:B::::::"),
	(0,     1,     0,     '*',     6,     0, ":::B::WW:B::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     0, "::::::::::B:::::"),
	(0,     0,     0,     'B',     0,     0, "::::::::::B:::::"),
	(0,     0,     1,     ':',     0,     0, "::::::::::B:::::"),
	(0,     0,     0,     '*',     15,     0, "::::::::::B:::::"),
	(0,     0,     0,     'W',     0,     0, "::::::::::B:::::"),
	(0,     1,     1,     ':',     10,     0, "::::::::::B:::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     3,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     2,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     7,     0, "::*:::::::::W:::"),
	(0,     0,     0,     ':',     0,     0, "::*::::*::::W:::"),
	(0,     0,     0,     'W',     12,     0, "::*::::*::::W:::"),
	(0,     1,     1,     'B',     0,     0, "::*::::*::::W:::"),
	(0,     0,     1,     '*',     10,     0, "B:::::::::::::::"),
	(0,     0,     0,     '*',     6,     0, "B:::::::::*:::::"),
	(0,     0,     0,     'B',     12,     0, "B:::::::::*:::::"),
	(0,     0,     0,     '*',     4,     0, "B:::::::::*:::::"),
	(0,     0,     0,     'W',     4,     0, "B:::::::::*:::::"),
	(0,     0,     1,     '*',     3,     0, "B:::::::::*:::::"),
	(0,     0,     1,     'W',     12,     0, "B::*::::::*:::::"),
	(0,     0,     0,     ':',     7,     0, "B::*::::::*:W:::"),
	(0,     0,     0,     ':',     7,     0, "B::*::::::*:W:::"),
	(0,     0,     0,     ':',     9,     0, "B::*::::::*:W:::"),
	(0,     0,     1,     ':',     5,     0, "B::*::::::*:W:::"),
	(0,     0,     1,     ':',     2,     0, "B::*::::::*:W:::"),
	(0,     0,     1,     'W',     5,     0, "B::*::::::*:W:::"),
	(0,     0,     0,     '*',     6,     0, "B::*:W::::*:W:::"),
	(0,     0,     0,     'B',     2,     0, "B::*:W::::*:W:::"),
	(0,     0,     1,     'W',     3,     0, "B::*:W::::*:W:::"),
	(0,     0,     1,     'B',     12,     0, "B::W:W::::*:W:::"),
	(0,     0,     1,     'W',     3,     0, "B::W:W::::*:B:::"),
	(0,     0,     0,     'W',     14,     0, "B::W:W::::*:B:::"),
	(0,     0,     0,     'B',     8,     0, "B::W:W::::*:B:::"),
	(0,     0,     1,     'W',     11,     0, "B::W:W::::*:B:::"),
	(0,     0,     0,     '*',     7,     0, "B::W:W::::*WB:::"),
	(0,     0,     0,     'W',     7,     0, "B::W:W::::*WB:::"),
	(0,     0,     1,     'W',     11,     0, "B::W:W::::*WB:::"),
	(0,     0,     0,     'B',     12,     0, "B::W:W::::*WB:::"),
	(0,     0,     0,     ':',     13,     0, "B::W:W::::*WB:::"),
	(0,     0,     1,     ':',     8,     0, "B::W:W::::*WB:::"),
	(0,     0,     1,     '*',     4,     0, "B::W:W::::*WB:::"),
	(0,     1,     1,     'W',     8,     0, "B::W*W::::*WB:::"),
	(0,     0,     1,     ':',     1,     0, "::::::::W:::::::"),
	(0,     0,     1,     'W',     10,     0, "::::::::W:::::::"),
	(0,     1,     1,     '*',     11,     0, "::::::::W:W:::::"),
	(0,     0,     0,     'B',     0,     0, ":::::::::::*::::"),
	(0,     1,     1,     'W',     10,     0, ":::::::::::*::::"),
	(0,     0,     0,     '*',     6,     0, "::::::::::W:::::"),
	(0,     0,     1,     'W',     5,     0, "::::::::::W:::::"),
	(0,     1,     1,     'W',     14,     0, ":::::W::::W:::::"),
	(0,     0,     1,     '*',     4,     0, "::::::::::::::W:"),
	(0,     0,     1,     'W',     15,     0, "::::*:::::::::W:"),
	(0,     0,     1,     ':',     13,     0, "::::*:::::::::WW"),
	(0,     0,     0,     'W',     12,     0, "::::*:::::::::WW"),
	(0,     0,     1,     '*',     9,     0, "::::*:::::::::WW"),
	(0,     0,     1,     'B',     5,     0, "::::*::::*::::WW"),
	(0,     0,     1,     'W',     11,     0, "::::*B:::*::::WW"),
	(0,     0,     0,     'B',     6,     0, "::::*B:::*:W::WW"),
	(0,     0,     0,     ':',     8,     0, "::::*B:::*:W::WW"),
	(0,     0,     1,     'W',     2,     0, "::::*B:::*:W::WW"),
	(0,     0,     1,     ':',     1,     0, "::W:*B:::*:W::WW"),
	(0,     0,     0,     'B',     3,     0, "::W:*B:::*:W::WW"),
	(0,     0,     0,     'B',     11,     0, "::W:*B:::*:W::WW"),
	(0,     0,     1,     '*',     14,     0, "::W:*B:::*:W::WW"),
	(0,     1,     1,     '*',     3,     0, "::W:*B:::*:W::BW"),
	(0,     0,     0,     'W',     12,     0, ":::*::::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     9,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     14,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::*::::::::::::"),
	(0,     0,     1,     '*',     6,     0, ":::*::::::::::::"),
	(0,     1,     0,     'B',     12,     0, ":::*::*:::::::::"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, ":::*::::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::*::::::::::::"),
	(0,     0,     0,     ':',     2,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     14,     0, ":::*::::::::::::"),
	(0,     0,     1,     'B',     4,     0, ":::*::::::::::::"),
	(0,     0,     1,     '*',     0,     0, ":::*B:::::::::::"),
	(0,     0,     1,     '*',     9,     0, "*::*B:::::::::::"),
	(0,     0,     1,     'B',     9,     0, "*::*B::::*::::::"),
	(0,     1,     1,     'W',     2,     0, "*::*B::::B::::::"),
	(0,     1,     0,     '*',     4,     0, "::W:::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     0, ":::::::::B::::::"),
	(0,     0,     1,     ':',     10,     0, ":::::::::B::::::"),
	(0,     0,     0,     ':',     12,     0, ":::::::::B::::::"),
	(0,     0,     0,     'B',     7,     0, ":::::::::B::::::"),
	(0,     1,     0,     'W',     10,     0, ":::::::::B::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     0, "::::::::::::B:::"),
	(0,     0,     1,     'B',     3,     0, "::::::::::::B:::"),
	(0,     0,     1,     ':',     13,     0, ":::B::::::::B:::"),
	(0,     0,     0,     '*',     3,     0, ":::B::::::::B:::"),
	(0,     0,     1,     ':',     0,     0, ":::B::::::::B:::"),
	(0,     0,     0,     ':',     6,     0, ":::B::::::::B:::"),
	(0,     0,     1,     'B',     10,     0, ":::B::::::::B:::"),
	(0,     0,     1,     '*',     2,     0, ":::B::::::B:B:::"),
	(0,     0,     1,     ':',     11,     0, "::*B::::::B:B:::"),
	(1,     0,     1,     ':',     9,     0, "::*B::::::B:B:::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     11,     0, ":::::*::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":::::*::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     8,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     7,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     2,     0, ":::::*::::::::::"),
	(0,     0,     0,     '*',     14,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     7,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::::*::::::::::"),
	(0,     0,     1,     ':',     10,     0, ":::::*::::::::::"),
	(0,     1,     1,     '*',     15,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::::::*"),
	(0,     0,     1,     '*',     0,     0, ":::::::::::::::*"),
	(0,     0,     1,     'W',     13,     0, "*::::::::::::::*"),
	(0,     0,     0,     ':',     0,     0, "*::::::::::::W:*"),
	(0,     0,     0,     'W',     5,     0, "*::::::::::::W:*"),
	(0,     0,     0,     ':',     15,     0, "*::::::::::::W:*"),
	(0,     0,     0,     'W',     12,     0, "*::::::::::::W:*"),
	(0,     0,     0,     ':',     13,     0, "*::::::::::::W:*"),
	(0,     0,     0,     ':',     1,     0, "*::::::::::::W:*"),
	(0,     0,     0,     'B',     1,     0, "*::::::::::::W:*"),
	(0,     0,     0,     'W',     8,     0, "*::::::::::::W:*"),
	(0,     0,     1,     ':',     14,     0, "*::::::::::::W:*"),
	(0,     0,     0,     ':',     5,     0, "*::::::::::::W:*"),
	(0,     0,     0,     'W',     11,     0, "*::::::::::::W:*"),
	(0,     0,     0,     ':',     15,     0, "*::::::::::::W:*"),
	(0,     0,     1,     'W',     9,     0, "*::::::::::::W:*"),
	(0,     0,     0,     'W',     14,     0, "*::::::::W:::W:*"),
	(0,     0,     1,     '*',     12,     0, "*::::::::W:::W:*"),
	(0,     0,     1,     'W',     2,     0, "*::::::::W::*W:*"),
	(0,     0,     0,     ':',     14,     0, "*:W::::::W::*W:*"),
	(0,     0,     0,     'B',     3,     0, "*:W::::::W::*W:*"),
	(0,     0,     0,     'B',     7,     0, "*:W::::::W::*W:*"),
	(0,     0,     0,     '*',     4,     0, "*:W::::::W::*W:*"),
	(0,     0,     1,     '*',     5,     0, "*:W::::::W::*W:*"),
	(0,     0,     1,     'W',     8,     0, "*:W::*:::W::*W:*"),
	(0,     0,     1,     'B',     9,     0, "*:W::*::WW::*W:*"),
	(0,     0,     1,     ':',     15,     0, "*:W::*::WB::*W:*"),
	(0,     0,     0,     'W',     11,     0, "*:W::*::WB::*W:*"),
	(0,     0,     1,     'W',     11,     0, "*:W::*::WB::*W:*"),
	(0,     1,     1,     'B',     0,     0, "*:W::*::WB:W*W:*"),
	(0,     0,     1,     'W',     7,     0, "B:::::::::::::::"),
	(0,     0,     0,     'W',     12,     0, "B::::::W::::::::"),
	(0,     0,     1,     'B',     9,     0, "B::::::W::::::::"),
	(0,     1,     0,     'B',     11,     0, "B::::::W:B::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     8,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     0, ":::W::::::::::::"),
	(0,     0,     1,     ':',     1,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::W::::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::W::::::::::::"),
	(0,     0,     1,     'B',     0,     0, ":::W::::::::::W:"),
	(0,     0,     1,     'W',     13,     0, "B::W::::::::::W:"),
	(1,     0,     1,     'B',     13,     0, "B::W:::::::::WW:"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, "*:::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "*::B::::::::::::"),
	(0,     0,     0,     '*',     5,     0, "*::B::::::::::::"),
	(0,     0,     1,     ':',     13,     0, "*::B::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "*::B::::::::::::"),
	(0,     0,     0,     'W',     3,     0, "*::B::::::::::::"),
	(0,     0,     1,     'B',     15,     0, "*::B::::::::::::"),
	(0,     0,     1,     ':',     14,     0, "*::B:::::::::::B"),
	(0,     0,     0,     'W',     8,     0, "*::B:::::::::::B"),
	(0,     0,     0,     'B',     4,     0, "*::B:::::::::::B"),
	(0,     0,     0,     '*',     10,     0, "*::B:::::::::::B"),
	(0,     0,     0,     ':',     6,     0, "*::B:::::::::::B"),
	(0,     0,     0,     '*',     7,     0, "*::B:::::::::::B"),
	(0,     0,     0,     ':',     8,     0, "*::B:::::::::::B"),
	(0,     0,     1,     'W',     13,     0, "*::B:::::::::::B"),
	(0,     0,     0,     '*',     0,     0, "*::B:::::::::W:B"),
	(0,     0,     1,     '*',     15,     0, "*::B:::::::::W:B"),
	(0,     0,     0,     ':',     8,     0, "*::B:::::::::W:W"),
	(0,     0,     0,     '*',     3,     0, "*::B:::::::::W:W"),
	(0,     0,     1,     ':',     1,     0, "*::B:::::::::W:W"),
	(0,     0,     0,     'W',     13,     0, "*::B:::::::::W:W"),
	(0,     0,     1,     ':',     6,     0, "*::B:::::::::W:W"),
	(0,     0,     0,     'W',     11,     0, "*::B:::::::::W:W"),
	(0,     0,     0,     'W',     14,     0, "*::B:::::::::W:W"),
	(0,     0,     0,     'W',     12,     0, "*::B:::::::::W:W"),
	(0,     0,     1,     '*',     13,     0, "*::B:::::::::W:W"),
	(0,     0,     0,     '*',     9,     0, "*::B:::::::::B:W"),
	(0,     0,     0,     '*',     14,     0, "*::B:::::::::B:W"),
	(0,     0,     1,     ':',     14,     0, "*::B:::::::::B:W"),
	(0,     0,     1,     'B',     1,     0, "*::B:::::::::B:W"),
	(0,     0,     0,     'W',     7,     0, "*B:B:::::::::B:W"),
	(0,     0,     0,     'B',     7,     0, "*B:B:::::::::B:W"),
	(0,     0,     0,     'B',     3,     0, "*B:B:::::::::B:W"),
	(0,     0,     1,     'W',     3,     0, "*B:B:::::::::B:W"),
	(0,     0,     0,     '*',     9,     0, "*B:W:::::::::B:W"),
	(0,     0,     0,     'B',     1,     0, "*B:W:::::::::B:W"),
	(0,     0,     1,     '*',     11,     0, "*B:W:::::::::B:W"),
	(0,     0,     1,     'B',     3,     0, "*B:W:::::::*:B:W"),
	(0,     0,     1,     'B',     14,     0, "*B:B:::::::*:B:W"),
	(0,     0,     1,     '*',     3,     0, "*B:B:::::::*:BBW"),
	(0,     0,     0,     'B',     6,     0, "*B:W:::::::*:BBW"),
	(0,     1,     0,     ':',     12,     0, "*B:W:::::::*:BBW"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     0, ":::::::::::W::::"),
	(0,     0,     1,     '*',     1,     0, ":::::::::B:W::::"),
	(0,     0,     0,     ':',     1,     0, ":*:::::::B:W::::"),
	(0,     0,     0,     ':',     1,     0, ":*:::::::B:W::::"),
	(0,     0,     0,     ':',     8,     0, ":*:::::::B:W::::"),
	(0,     1,     1,     ':',     8,     0, ":*:::::::B:W::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, "::W:::::::::::::"),
	(0,     0,     1,     'B',     7,     0, "::W:::::::::::::"),
	(0,     0,     1,     'W',     5,     0, "::W::::B::::::::"),
	(0,     0,     0,     '*',     12,     0, "::W::W:B::::::::"),
	(0,     0,     0,     'W',     2,     0, "::W::W:B::::::::"),
	(0,     0,     0,     'B',     4,     0, "::W::W:B::::::::"),
	(0,     1,     0,     '*',     8,     0, "::W::W:B::::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     0, ":::::::B::::::::"),
	(0,     0,     0,     '*',     11,     0, ":::::::B::::::::"),
	(0,     0,     1,     'W',     12,     0, ":::::::B::::::::"),
	(0,     0,     1,     '*',     9,     0, ":::::::B::::W:::"),
	(0,     0,     1,     ':',     11,     0, ":::::::B:*::W:::"),
	(0,     1,     1,     '*',     2,     0, ":::::::B:*::W:::"),
	(0,     0,     1,     'B',     3,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "::*B::::::::::::"),
	(1,     0,     0,     'W',     10,     0, "::*B::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     12,     0, "::::::::::::::B:"),
	(0,     0,     1,     'B',     9,     0, "::::::::::::W:B:"),
	(0,     1,     1,     ':',     14,     0, ":::::::::B::W:B:"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     0, ":::::*::::::::::"),
	(0,     0,     0,     '*',     15,     0, ":::::*::::::::::"),
	(0,     1,     0,     '*',     10,     0, ":::::*::::::::::"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     5,     0, ":::B::::::::::::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     0, ":::::::::*::::::"),
	(0,     0,     1,     'B',     13,     0, ":::::::::*::::::"),
	(0,     0,     1,     'W',     9,     0, ":::::::::*:::B::"),
	(0,     1,     0,     '*',     11,     0, ":::::::::W:::B::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     12,     0, ":::::B::::::::::"),
	(0,     0,     0,     ':',     14,     0, ":::::B::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::::B::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::::B::::::::::"),
	(0,     0,     0,     'W',     0,     0, ":::::B::::::::W:"),
	(0,     0,     0,     'B',     10,     0, ":::::B::::::::W:"),
	(0,     0,     0,     'B',     15,     0, ":::::B::::::::W:"),
	(0,     0,     1,     ':',     5,     0, ":::::B::::::::W:"),
	(0,     0,     0,     ':',     8,     0, ":::::B::::::::W:"),
	(0,     0,     1,     '*',     7,     0, ":::::B::::::::W:"),
	(0,     0,     1,     'B',     11,     0, ":::::B:*::::::W:"),
	(0,     0,     0,     'W',     4,     0, ":::::B:*:::B::W:"),
	(0,     0,     0,     ':',     1,     0, ":::::B:*:::B::W:"),
	(0,     0,     1,     '*',     1,     0, ":::::B:*:::B::W:"),
	(0,     0,     1,     ':',     1,     0, ":*:::B:*:::B::W:"),
	(0,     0,     0,     'B',     5,     0, ":*:::B:*:::B::W:"),
	(0,     0,     1,     'W',     10,     0, ":*:::B:*:::B::W:"),
	(0,     0,     0,     'W',     7,     0, ":*:::B:*::WB::W:"),
	(0,     0,     0,     'B',     2,     0, ":*:::B:*::WB::W:"),
	(0,     0,     1,     '*',     7,     0, ":*:::B:*::WB::W:"),
	(0,     0,     0,     '*',     11,     0, ":*:::B::::WB::W:"),
	(0,     0,     1,     '*',     6,     0, ":*:::B::::WB::W:"),
	(0,     0,     0,     '*',     10,     0, ":*:::B*:::WB::W:"),
	(0,     0,     1,     '*',     0,     0, ":*:::B*:::WB::W:"),
	(0,     1,     0,     ':',     9,     0, "**:::B*:::WB::W:"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     1,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     12,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::*:::::::::B:::"),
	(0,     0,     0,     'B',     15,     0, "::*:::::::::B:::"),
	(0,     0,     1,     'B',     3,     0, "::*:::::::::B:::"),
	(0,     1,     0,     '*',     7,     0, "::*B::::::::B:::"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, ":::::::B::::::::"),
	(0,     0,     0,     '*',     4,     0, ":::::::B::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::::::B::::::::"),
	(0,     1,     0,     ':',     15,     0, ":::::::B::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     0, "*:::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "*::::::::W::::::"),
	(0,     0,     0,     'W',     3,     0, "*::::::::W::::::"),
	(0,     0,     1,     ':',     8,     0, "*::::::::W::::::"),
	(0,     1,     0,     'B',     4,     0, "*::::::::W::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     0, "::::::::::::::W:"),
	(0,     0,     1,     ':',     4,     0, "::::::::::::::W:"),
	(0,     0,     0,     '*',     0,     0, "::::::::::::::W:"),
	(0,     0,     1,     'B',     0,     0, "::::::::::::::W:"),
	(0,     0,     0,     'W',     12,     0, "B:::::::::::::W:"),
	(0,     0,     1,     'B',     15,     0, "B:::::::::::::W:"),
	(0,     0,     0,     '*',     14,     0, "B:::::::::::::WB"),
	(0,     0,     1,     '*',     5,     0, "B:::::::::::::WB"),
	(0,     0,     1,     'B',     2,     0, "B::::*::::::::WB"),
	(0,     0,     0,     'W',     13,     0, "B:B::*::::::::WB"),
	(0,     0,     0,     '*',     0,     0, "B:B::*::::::::WB"),
	(0,     0,     1,     '*',     4,     0, "B:B::*::::::::WB"),
	(0,     1,     0,     'B',     9,     0, "B:B:**::::::::WB"),
	(0,     1,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     1,     0, "::B:::B:::::::::"),
	(0,     0,     1,     'B',     9,     0, "::B:::B:::::::::"),
	(0,     1,     1,     'B',     13,     0, "::B:::B::B::::::"),
	(0,     0,     0,     ':',     11,     0, ":::::::::::::B::"),
	(0,     0,     0,     ':',     9,     0, ":::::::::::::B::"),
	(0,     0,     0,     '*',     4,     0, ":::::::::::::B::"),
	(0,     0,     0,     'B',     7,     0, ":::::::::::::B::"),
	(0,     0,     0,     '*',     2,     0, ":::::::::::::B::"),
	(0,     0,     0,     'B',     7,     0, ":::::::::::::B::"),
	(0,     0,     1,     '*',     12,     0, ":::::::::::::B::"),
	(0,     0,     1,     '*',     10,     0, "::::::::::::*B::"),
	(0,     0,     0,     'W',     2,     0, "::::::::::*:*B::"),
	(0,     0,     1,     '*',     11,     0, "::::::::::*:*B::"),
	(0,     0,     0,     ':',     15,     0, "::::::::::***B::"),
	(0,     0,     0,     '*',     4,     0, "::::::::::***B::"),
	(0,     0,     1,     ':',     3,     0, "::::::::::***B::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::***B::"),
	(0,     0,     0,     '*',     5,     0, "::::::::::***B::"),
	(0,     0,     0,     '*',     0,     0, "::::::::::***B::"),
	(0,     0,     1,     '*',     9,     0, "::::::::::***B::"),
	(0,     0,     1,     '*',     13,     0, ":::::::::****B::"),
	(0,     0,     0,     'B',     6,     0, ":::::::::****W::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::****W::"),
	(0,     0,     1,     '*',     12,     0, "::::::::*****W::"),
	(0,     0,     0,     'W',     0,     0, "::::::::****:W::"),
	(0,     0,     0,     'B',     4,     0, "::::::::****:W::"),
	(0,     0,     0,     'B',     10,     0, "::::::::****:W::"),
	(0,     0,     0,     '*',     10,     0, "::::::::****:W::"),
	(0,     0,     0,     'B',     3,     0, "::::::::****:W::"),
	(0,     0,     1,     'B',     9,     0, "::::::::****:W::"),
	(0,     0,     1,     ':',     9,     0, "::::::::*B**:W::"),
	(0,     0,     1,     '*',     8,     0, "::::::::*B**:W::"),
	(0,     1,     0,     '*',     11,     0, ":::::::::B**:W::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     0, "::::::::::::B:::"),
	(0,     0,     0,     'B',     2,     0, "::::::::::::B:::"),
	(0,     1,     0,     '*',     10,     0, "::::::::::::B:::"),
	(0,     0,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::B:::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::B:::::::::"),
	(0,     0,     0,     ':',     13,     0, "::::::B:::::::::"),
	(0,     0,     1,     '*',     13,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     3,     0, "::::::B::::::*::"),
	(0,     0,     1,     '*',     12,     0, "::::::B::::::*::"),
	(0,     0,     1,     ':',     11,     0, "::::::B:::::**::"),
	(0,     1,     0,     'B',     5,     0, "::::::B:::::**::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     12,     0, ":::::::*::::::::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::::B:::"),
	(0,     0,     0,     '*',     15,     0, "::::::::::::B:::"),
	(0,     0,     1,     ':',     4,     0, "::::::::::::B:::"),
	(0,     0,     0,     'B',     4,     0, "::::::::::::B:::"),
	(0,     0,     0,     ':',     10,     0, "::::::::::::B:::"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::B:::"),
	(0,     0,     0,     'W',     2,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     12,     0, "::::::::::::B:::"),
	(0,     0,     0,     ':',     15,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     5,     0, "::::::::::::W:::"),
	(1,     0,     0,     'W',     3,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(1,     1,     0,     'B',     5,     1, "::::::::::::::::"),
	(1,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, ":::::B::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::::B::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     14,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":::::B::::::::B:"),
	(0,     0,     1,     ':',     1,     0, ":::::B:::::::*B:"),
	(0,     0,     1,     'B',     7,     0, ":::::B:::::::*B:"),
	(0,     0,     0,     'B',     4,     0, ":::::B:B:::::*B:"),
	(0,     0,     0,     'B',     15,     0, ":::::B:B:::::*B:"),
	(0,     1,     0,     ':',     1,     0, ":::::B:B:::::*B:"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::::W::::::::W:"),
	(0,     0,     0,     ':',     6,     0, ":::::W::::::::W:"),
	(0,     0,     0,     ':',     6,     0, ":::::W::::::::W:"),
	(0,     0,     1,     'W',     5,     0, ":::::W::::::::W:"),
	(0,     0,     0,     ':',     8,     0, ":::::W::::::::W:"),
	(0,     0,     1,     '*',     15,     0, ":::::W::::::::W:"),
	(0,     1,     1,     ':',     9,     0, ":::::W::::::::W*"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     0,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     9,     0, "W:::::::::::B:::"),
	(0,     1,     0,     ':',     7,     0, "W::::::::W::B:::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     0, "W:::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "W:::B:::::::::::"),
	(0,     0,     0,     'W',     12,     0, "W:::B:::::::::::"),
	(0,     0,     1,     'B',     7,     0, "W:::B:::::::::::"),
	(0,     0,     0,     'B',     12,     0, "W:::B::B::::::::"),
	(0,     0,     0,     'W',     5,     0, "W:::B::B::::::::"),
	(0,     0,     1,     'W',     9,     0, "W:::B::B::::::::"),
	(0,     0,     1,     'W',     9,     0, "W:::B::B:W::::::"),
	(0,     0,     1,     'B',     14,     0, "W:::B::B:W::::::"),
	(0,     0,     0,     'W',     11,     0, "W:::B::B:W::::B:"),
	(0,     0,     1,     ':',     9,     0, "W:::B::B:W::::B:"),
	(0,     0,     1,     '*',     5,     0, "W:::B::B:W::::B:"),
	(0,     0,     1,     '*',     4,     0, "W:::B*:B:W::::B:"),
	(0,     0,     0,     'W',     8,     0, "W:::W*:B:W::::B:"),
	(0,     0,     1,     ':',     10,     0, "W:::W*:B:W::::B:"),
	(0,     0,     0,     ':',     14,     0, "W:::W*:B:W::::B:"),
	(0,     0,     1,     'B',     10,     0, "W:::W*:B:W::::B:"),
	(0,     0,     1,     'W',     13,     0, "W:::W*:B:WB:::B:"),
	(0,     0,     0,     ':',     8,     0, "W:::W*:B:WB::WB:"),
	(0,     0,     0,     '*',     13,     0, "W:::W*:B:WB::WB:"),
	(0,     0,     0,     'B',     8,     0, "W:::W*:B:WB::WB:"),
	(0,     1,     0,     '*',     7,     0, "W:::W*:B:WB::WB:"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     10,     0, "::::::::::W:::::"),
	(0,     0,     1,     'W',     12,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     11,     0, "::::::::::W:W:::"),
	(0,     0,     1,     'W',     6,     0, "::::::::::W:W:::"),
	(0,     0,     1,     'W',     13,     0, "::::::W:::W:W:::"),
	(0,     0,     0,     'W',     3,     0, "::::::W:::W:WW::"),
	(0,     0,     0,     'W',     6,     0, "::::::W:::W:WW::"),
	(0,     0,     0,     'W',     2,     0, "::::::W:::W:WW::"),
	(0,     0,     1,     'B',     11,     0, "::::::W:::W:WW::"),
	(0,     0,     0,     '*',     2,     0, "::::::W:::WBWW::"),
	(0,     0,     1,     '*',     5,     0, "::::::W:::WBWW::"),
	(0,     1,     0,     'B',     13,     0, ":::::*W:::WBWW::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, ":B::::::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":B::::::B:::::::"),
	(0,     0,     0,     'B',     5,     0, ":B::::::B:::::::"),
	(0,     1,     1,     'W',     8,     0, ":B::::::B:::::::"),
	(0,     0,     0,     'W',     6,     0, "::::::::W:::::::"),
	(0,     1,     0,     ':',     4,     0, "::::::::W:::::::"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     13,     0, "::::::::::::B:::"),
	(0,     0,     0,     '*',     6,     0, "::::::::::::BW::"),
	(0,     0,     0,     'W',     2,     0, "::::::::::::BW::"),
	(0,     0,     1,     'B',     6,     0, "::::::::::::BW::"),
	(0,     0,     0,     'W',     10,     0, "::::::B:::::BW::"),
	(0,     0,     1,     'W',     11,     0, "::::::B:::::BW::"),
	(0,     0,     1,     '*',     4,     0, "::::::B::::WBW::"),
	(0,     0,     0,     ':',     15,     0, "::::*:B::::WBW::"),
	(0,     0,     0,     'W',     2,     0, "::::*:B::::WBW::"),
	(0,     0,     1,     'B',     2,     0, "::::*:B::::WBW::"),
	(0,     0,     0,     '*',     5,     0, "::B:*:B::::WBW::"),
	(0,     0,     0,     '*',     0,     0, "::B:*:B::::WBW::"),
	(0,     0,     0,     'W',     1,     0, "::B:*:B::::WBW::"),
	(0,     1,     0,     'W',     4,     0, "::B:*:B::::WBW::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     0, ":::W::::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":::W::::::::::::"),
	(0,     0,     0,     '*',     1,     0, ":::W::::::::*:::"),
	(0,     0,     0,     '*',     11,     0, ":::W::::::::*:::"),
	(0,     0,     1,     '*',     4,     0, ":::W::::::::*:::"),
	(0,     0,     0,     'W',     10,     0, ":::W*:::::::*:::"),
	(0,     0,     1,     '*',     15,     0, ":::W*:::::::*:::"),
	(0,     0,     0,     '*',     0,     0, ":::W*:::::::*::*"),
	(0,     1,     1,     ':',     14,     0, ":::W*:::::::*::*"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     0, ":::::B::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::B::::::::::"),
	(0,     0,     0,     '*',     3,     0, ":::::B::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::::B::::::::::"),
	(0,     0,     1,     ':',     3,     0, ":::::B:::::::::W"),
	(0,     0,     0,     '*',     2,     0, ":::::B:::::::::W"),
	(0,     0,     0,     '*',     13,     0, ":::::B:::::::::W"),
	(0,     0,     0,     ':',     8,     0, ":::::B:::::::::W"),
	(0,     0,     1,     '*',     7,     0, ":::::B:::::::::W"),
	(0,     0,     1,     'B',     9,     0, ":::::B:*:::::::W"),
	(0,     0,     0,     'B',     12,     0, ":::::B:*:B:::::W"),
	(0,     0,     0,     ':',     12,     0, ":::::B:*:B:::::W"),
	(0,     0,     0,     '*',     7,     0, ":::::B:*:B:::::W"),
	(0,     0,     0,     ':',     3,     0, ":::::B:*:B:::::W"),
	(0,     0,     0,     'W',     5,     0, ":::::B:*:B:::::W"),
	(0,     1,     1,     'B',     10,     0, ":::::B:*:B:::::W"),
	(0,     0,     0,     'W',     10,     0, "::::::::::B:::::"),
	(0,     0,     1,     'W',     5,     0, "::::::::::B:::::"),
	(0,     1,     0,     'B',     2,     0, ":::::W::::B:::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     0, ":::::::::::::W::"),
	(0,     1,     1,     'W',     9,     0, ":::::::::::::W::"),
	(0,     0,     0,     ':',     15,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     14,     0, ":::::::::W::::::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::W::::::"),
	(0,     0,     0,     'B',     5,     0, ":::::::::W::::::"),
	(0,     0,     0,     '*',     5,     0, ":::::::::W::::::"),
	(0,     0,     1,     'W',     3,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     13,     0, ":::W:::::W::::::"),
	(0,     0,     1,     ':',     12,     0, ":::W:::::W::::::"),
	(0,     0,     0,     'B',     9,     0, ":::W:::::W::::::"),
	(0,     0,     0,     ':',     15,     0, ":::W:::::W::::::"),
	(0,     1,     0,     'W',     1,     0, ":::W:::::W::::::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     11,     0, "::::::::::::*:::"),
	(0,     0,     0,     ':',     0,     0, "::::::::::::*:::"),
	(0,     0,     0,     'W',     6,     0, "::::::::::::*:::"),
	(0,     0,     1,     '*',     0,     0, "::::::::::::*:::"),
	(0,     1,     0,     ':',     1,     0, "*:::::::::::*:::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::::::W:::::::::"),
	(0,     0,     0,     '*',     11,     0, "::::::W:::::::W:"),
	(0,     0,     1,     '*',     12,     0, "::::::W:::::::W:"),
	(0,     0,     1,     ':',     10,     0, "::::::W:::::*:W:"),
	(0,     0,     0,     '*',     7,     0, "::::::W:::::*:W:"),
	(0,     0,     1,     'B',     14,     0, "::::::W:::::*:W:"),
	(0,     0,     1,     '*',     2,     0, "::::::W:::::*:B:"),
	(0,     0,     1,     'B',     12,     0, "::*:::W:::::*:B:"),
	(0,     0,     1,     ':',     0,     0, "::*:::W:::::B:B:"),
	(0,     0,     1,     '*',     6,     0, "::*:::W:::::B:B:"),
	(0,     0,     0,     '*',     11,     0, "::*:::B:::::B:B:"),
	(0,     0,     0,     ':',     3,     0, "::*:::B:::::B:B:"),
	(0,     0,     1,     '*',     4,     0, "::*:::B:::::B:B:"),
	(0,     0,     1,     'W',     10,     0, "::*:*:B:::::B:B:"),
	(0,     1,     0,     ':',     2,     0, "::*:*:B:::W:B:B:"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     1,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     9,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     11,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     6,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     11,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, "*:::::::::::::::"),
	(0,     0,     0,     ':',     14,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     7,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     4,     0, "*:::::::::::::::"),
	(0,     0,     0,     ':',     6,     0, "*:::::::::::::::"),
	(0,     1,     0,     'W',     6,     0, "*:::::::::::::::"),
	(0,     0,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::::::::::::::*"),
	(0,     1,     0,     'B',     6,     0, ":::::::::::::::*"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     3,     0, ":::::::::*::::::"),
	(0,     0,     0,     ':',     12,     0, ":::*:::::*::::::"),
	(0,     1,     0,     'B',     4,     0, ":::*:::::*::::::"),
	(0,     1,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     0, "::::::::::::::W:"),
	(0,     0,     1,     ':',     1,     0, "::::::::::::W:W:"),
	(0,     1,     1,     'W',     2,     0, "::::::::::::W:W:"),
	(0,     0,     1,     'W',     10,     0, "::W:::::::::::::"),
	(0,     0,     0,     ':',     14,     0, "::W:::::::W:::::"),
	(0,     0,     0,     ':',     15,     0, "::W:::::::W:::::"),
	(0,     1,     1,     ':',     9,     0, "::W:::::::W:::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     0, "W:::::::::::::::"),
	(0,     0,     1,     ':',     12,     0, "W:::::::::::::::"),
	(0,     0,     0,     'W',     5,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     5,     0, "W:::::::::::::::"),
	(0,     1,     0,     'B',     3,     0, "W::::*::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     15,     0, ":::::::::::::::W"),
	(0,     0,     1,     'W',     12,     0, ":::::::::::::::B"),
	(0,     0,     1,     'W',     5,     0, "::::::::::::W::B"),
	(0,     1,     0,     ':',     6,     0, ":::::W::::::W::B"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, "::::::W:::::::::"),
	(0,     0,     1,     '*',     4,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     12,     0, "::::*:W:::::::::"),
	(0,     0,     0,     'W',     8,     0, "::::*:W:::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::*:W:::::::::"),
	(0,     0,     1,     ':',     9,     0, "::*:*:W:::::::::"),
	(0,     0,     0,     ':',     12,     0, "::*:*:W:::::::::"),
	(0,     0,     1,     'W',     10,     0, "::*:*:W:::::::::"),
	(0,     0,     0,     ':',     7,     0, "::*:*:W:::W:::::"),
	(0,     0,     0,     ':',     2,     0, "::*:*:W:::W:::::"),
	(0,     0,     1,     'W',     5,     0, "::*:*:W:::W:::::"),
	(0,     0,     1,     '*',     9,     0, "::*:*WW:::W:::::"),
	(0,     0,     0,     'B',     6,     0, "::*:*WW::*W:::::"),
	(0,     0,     0,     'B',     2,     0, "::*:*WW::*W:::::"),
	(0,     0,     0,     ':',     12,     0, "::*:*WW::*W:::::"),
	(0,     1,     0,     'W',     14,     0, "::*:*WW::*W:::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     0, ":::::::::::B::::"),
	(0,     0,     1,     ':',     12,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     0,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     14,     0, "*::::::::::B::::"),
	(0,     0,     0,     'B',     4,     0, "*::::::::::B::::"),
	(0,     0,     1,     'B',     9,     0, "*::::::::::B::::"),
	(0,     0,     1,     '*',     1,     0, "*::::::::B:B::::"),
	(0,     0,     1,     'W',     10,     0, "**:::::::B:B::::"),
	(0,     0,     0,     'B',     10,     0, "**:::::::BWB::::"),
	(0,     0,     0,     ':',     1,     0, "**:::::::BWB::::"),
	(0,     0,     1,     'B',     4,     0, "**:::::::BWB::::"),
	(0,     0,     0,     ':',     10,     0, "**::B::::BWB::::"),
	(1,     0,     1,     'B',     10,     0, "**::B::::BWB::::"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     12,     0, ":W::::::::::::::"),
	(0,     0,     1,     ':',     3,     0, "::::::::::::B:::"),
	(0,     0,     0,     'B',     1,     0, "::::::::::::B:::"),
	(0,     0,     1,     'B',     6,     0, "::::::::::::B:::"),
	(0,     0,     1,     ':',     2,     0, "::::::B:::::B:::"),
	(0,     1,     1,     'B',     7,     0, "::::::B:::::B:::"),
	(0,     0,     0,     'W',     9,     0, ":::::::B::::::::"),
	(0,     0,     1,     ':',     15,     0, ":::::::B::::::::"),
	(0,     0,     1,     '*',     4,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     1,     0, "::::*::B::::::::"),
	(0,     0,     1,     'W',     2,     0, "::::*::B::::::::"),
	(0,     0,     1,     'W',     13,     0, "::W:*::B::::::::"),
	(0,     0,     1,     'B',     12,     0, "::W:*::B:::::W::"),
	(0,     0,     0,     ':',     14,     0, "::W:*::B::::BW::"),
	(0,     0,     1,     ':',     4,     0, "::W:*::B::::BW::"),
	(0,     0,     0,     ':',     9,     0, "::W:*::B::::BW::"),
	(0,     0,     0,     'B',     11,     0, "::W:*::B::::BW::"),
	(0,     0,     0,     'W',     11,     0, "::W:*::B::::BW::"),
	(0,     1,     0,     'B',     2,     0, "::W:*::B::::BW::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     3,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     6,     0, ":::::::::::::::B"),
	(0,     0,     0,     ':',     12,     0, ":::::::::::::::B"),
	(0,     0,     1,     'B',     10,     0, ":::::::::::::::B"),
	(0,     0,     1,     'W',     11,     0, "::::::::::B::::B"),
	(0,     0,     1,     '*',     6,     0, "::::::::::BW:::B"),
	(0,     0,     0,     ':',     0,     0, "::::::*:::BW:::B"),
	(0,     0,     0,     '*',     3,     0, "::::::*:::BW:::B"),
	(0,     0,     1,     'W',     2,     0, "::::::*:::BW:::B"),
	(0,     0,     0,     'W',     0,     0, "::W:::*:::BW:::B"),
	(0,     0,     1,     'B',     11,     0, "::W:::*:::BW:::B"),
	(0,     1,     1,     '*',     15,     0, "::W:::*:::BB:::B"),
	(0,     0,     1,     ':',     12,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     5,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     11,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     12,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     12,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     1,     0, ":::::::::::::::*"),
	(0,     0,     1,     '*',     9,     0, ":::::::::::::::*"),
	(0,     0,     0,     'W',     2,     0, ":::::::::*:::::*"),
	(0,     0,     1,     'B',     10,     0, ":::::::::*:::::*"),
	(0,     0,     1,     'W',     11,     0, ":::::::::*B::::*"),
	(0,     0,     1,     'B',     13,     0, ":::::::::*BW:::*"),
	(0,     1,     1,     'B',     1,     0, ":::::::::*BW:B:*"),
	(0,     1,     0,     'W',     4,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, ":::::::::::::::*"),
	(0,     0,     1,     '*',     9,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     15,     0, ":::::::::*:::::*"),
	(0,     1,     1,     ':',     2,     0, ":::::::::*:::::*"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, ":::::::::::::W::"),
	(0,     0,     1,     '*',     2,     0, ":::::::::::::W::"),
	(0,     0,     1,     ':',     15,     0, "::*::::::::::W::"),
	(0,     0,     1,     ':',     1,     0, "::*::::::::::W::"),
	(0,     0,     1,     'B',     9,     0, "::*::::::::::W::"),
	(0,     0,     1,     'W',     4,     0, "::*::::::B:::W::"),
	(0,     0,     0,     '*',     9,     0, "::*:W::::B:::W::"),
	(0,     0,     1,     'W',     3,     0, "::*:W::::B:::W::"),
	(0,     1,     0,     '*',     5,     0, "::*WW::::B:::W::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::::::W:::::::::"),
	(0,     0,     1,     '*',     15,     0, "::::::W:::::::W:"),
	(0,     0,     0,     '*',     6,     0, "::::::W:::::::W*"),
	(0,     0,     1,     ':',     1,     0, "::::::W:::::::W*"),
	(0,     0,     0,     '*',     15,     0, "::::::W:::::::W*"),
	(0,     0,     0,     'W',     3,     0, "::::::W:::::::W*"),
	(0,     0,     1,     '*',     7,     0, "::::::W:::::::W*"),
	(0,     0,     0,     'B',     0,     0, "::::::W*::::::W*"),
	(0,     1,     1,     'W',     13,     0, "::::::W*::::::W*"),
	(0,     0,     1,     'B',     9,     0, ":::::::::::::W::"),
	(0,     0,     1,     '*',     3,     0, ":::::::::B:::W::"),
	(0,     0,     0,     'B',     0,     0, ":::*:::::B:::W::"),
	(0,     0,     1,     ':',     1,     0, ":::*:::::B:::W::"),
	(0,     0,     1,     '*',     3,     0, ":::*:::::B:::W::"),
	(0,     0,     1,     '*',     5,     0, ":::::::::B:::W::"),
	(0,     0,     1,     '*',     7,     0, ":::::*:::B:::W::"),
	(0,     0,     0,     '*',     11,     0, ":::::*:*:B:::W::"),
	(0,     0,     0,     'B',     14,     0, ":::::*:*:B:::W::"),
	(0,     1,     1,     ':',     3,     0, ":::::*:*:B:::W::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::::::::::::*:::"),
	(0,     0,     1,     '*',     8,     0, "::::::::::::*:::"),
	(0,     0,     1,     'B',     7,     0, "::::::::*:::*:::"),
	(0,     1,     0,     'W',     2,     0, ":::::::B*:::*:::"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, "::W:::::::::::::"),
	(0,     0,     1,     ':',     11,     0, "::W:::::::::::::"),
	(0,     0,     1,     'B',     2,     0, "::W:::::::::::::"),
	(0,     1,     1,     'B',     14,     0, "::B:::::::::::::"),
	(0,     0,     1,     'B',     6,     0, "::::::::::::::B:"),
	(0,     1,     0,     'B',     13,     0, "::::::B:::::::B:"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     0, "B:::::::::::::::"),
	(0,     1,     0,     '*',     8,     0, "B:::::::::W:::::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     0,     0, "::::::::::::B:::"),
	(0,     0,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     13,     0, "::::::B:::::::::"),
	(0,     0,     0,     '*',     4,     0, "::::::B:::::::::"),
	(0,     0,     1,     '*',     0,     0, "::::::B:::::::::"),
	(0,     0,     1,     'W',     10,     0, "*:::::B:::::::::"),
	(0,     0,     1,     ':',     2,     0, "*:::::B:::W:::::"),
	(0,     0,     0,     'B',     6,     0, "*:::::B:::W:::::"),
	(0,     0,     1,     'B',     12,     0, "*:::::B:::W:::::"),
	(0,     0,     0,     'W',     15,     0, "*:::::B:::W:B:::"),
	(0,     0,     1,     'B',     13,     0, "*:::::B:::W:B:::"),
	(0,     0,     1,     '*',     5,     0, "*:::::B:::W:BB::"),
	(0,     0,     1,     ':',     15,     0, "*::::*B:::W:BB::"),
	(0,     0,     1,     ':',     4,     0, "*::::*B:::W:BB::"),
	(0,     0,     0,     '*',     8,     0, "*::::*B:::W:BB::"),
	(0,     0,     1,     'W',     12,     0, "*::::*B:::W:BB::"),
	(0,     1,     1,     '*',     12,     0, "*::::*B:::W:WB::"),
	(0,     1,     0,     '*',     10,     0, "::::::::::::*:::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     14,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":*::::::::::::B:"),
	(0,     0,     0,     '*',     8,     0, ":*::::::::::::B:"),
	(0,     0,     0,     ':',     15,     0, ":*::::::::::::B:"),
	(0,     0,     1,     '*',     4,     0, ":*::::::::::::B:"),
	(0,     0,     1,     '*',     6,     0, ":*::*:::::::::B:"),
	(0,     1,     1,     'W',     10,     0, ":*::*:*:::::::B:"),
	(0,     0,     0,     'W',     9,     0, "::::::::::W:::::"),
	(0,     0,     1,     'B',     3,     0, "::::::::::W:::::"),
	(0,     0,     0,     ':',     1,     0, ":::B::::::W:::::"),
	(0,     0,     0,     'W',     2,     0, ":::B::::::W:::::"),
	(0,     0,     0,     '*',     4,     0, ":::B::::::W:::::"),
	(0,     0,     1,     'B',     12,     0, ":::B::::::W:::::"),
	(0,     0,     1,     'B',     15,     0, ":::B::::::W:B:::"),
	(0,     1,     0,     'W',     1,     0, ":::B::::::W:B::B"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     2,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     11,     0, "::W::*::::::::::"),
	(0,     0,     0,     'B',     12,     0, "::W::*::::::::::"),
	(0,     0,     1,     'W',     8,     0, "::W::*::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::W::*::W:::::::"),
	(0,     1,     0,     ':',     12,     0, "::W::*::W:::::::"),
	(0,     0,     1,     '*',     13,     1, "::::::::::::::::"),
	(1,     1,     0,     'W',     4,     0, ":::::::::::::*::"),
	(0,     1,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::::::::::B::::"),
	(0,     0,     1,     ':',     1,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     1,     0, ":::::::::::B::::"),
	(0,     1,     1,     'W',     3,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     5,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     12,     0, ":::W:*::::::::::"),
	(0,     0,     0,     'W',     5,     0, ":::W:*::::::::::"),
	(0,     0,     0,     ':',     10,     0, ":::W:*::::::::::"),
	(0,     0,     0,     'W',     13,     0, ":::W:*::::::::::"),
	(0,     0,     0,     '*',     1,     0, ":::W:*::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::W:*::::::::::"),
	(0,     0,     1,     'W',     9,     0, ":::W:*::::::::::"),
	(0,     0,     1,     '*',     6,     0, ":::W:*:::W::::::"),
	(0,     0,     0,     '*',     8,     0, ":::W:**::W::::::"),
	(0,     0,     0,     'B',     7,     0, ":::W:**::W::::::"),
	(0,     0,     1,     ':',     15,     0, ":::W:**::W::::::"),
	(0,     0,     0,     ':',     14,     0, ":::W:**::W::::::"),
	(0,     1,     1,     'W',     15,     0, ":::W:**::W::::::"),
	(0,     0,     0,     'B',     9,     0, ":::::::::::::::W"),
	(0,     0,     1,     'W',     1,     0, ":::::::::::::::W"),
	(0,     0,     1,     '*',     1,     0, ":W:::::::::::::W"),
	(0,     0,     1,     'B',     10,     0, ":B:::::::::::::W"),
	(0,     0,     1,     'W',     14,     0, ":B::::::::B::::W"),
	(0,     0,     0,     'W',     14,     0, ":B::::::::B:::WW"),
	(0,     0,     0,     'B',     3,     0, ":B::::::::B:::WW"),
	(0,     0,     0,     'W',     6,     0, ":B::::::::B:::WW"),
	(0,     0,     0,     '*',     1,     0, ":B::::::::B:::WW"),
	(0,     0,     1,     'B',     0,     0, ":B::::::::B:::WW"),
	(0,     0,     0,     'B',     8,     0, "BB::::::::B:::WW"),
	(0,     0,     1,     'B',     8,     0, "BB::::::::B:::WW"),
	(0,     0,     0,     ':',     11,     0, "BB::::::B:B:::WW"),
	(0,     0,     1,     'W',     9,     0, "BB::::::B:B:::WW"),
	(0,     0,     1,     ':',     8,     0, "BB::::::BWB:::WW"),
	(0,     1,     1,     '*',     15,     0, "BB::::::BWB:::WW"),
	(0,     0,     0,     'B',     14,     0, ":::::::::::::::*"),
	(0,     1,     0,     'B',     12,     0, ":::::::::::::::*"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     10,     0, "B:::::::::::::B:"),
	(0,     1,     0,     'W',     0,     0, "B:::::::::::::B:"),
	(0,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     0,     0, "::::::::::::*:::"),
	(0,     0,     0,     'W',     11,     0, "::::::::::::*:::"),
	(0,     0,     1,     ':',     2,     0, "::::::::::::*:::"),
	(0,     0,     1,     'B',     9,     0, "::::::::::::*:::"),
	(0,     0,     1,     'W',     15,     0, ":::::::::B::*:::"),
	(0,     0,     1,     '*',     14,     0, ":::::::::B::*::W"),
	(0,     0,     0,     ':',     10,     0, ":::::::::B::*:*W"),
	(0,     0,     0,     '*',     11,     0, ":::::::::B::*:*W"),
	(0,     0,     0,     '*',     1,     0, ":::::::::B::*:*W"),
	(0,     0,     0,     'B',     6,     0, ":::::::::B::*:*W"),
	(0,     0,     0,     '*',     7,     0, ":::::::::B::*:*W"),
	(0,     0,     0,     ':',     0,     0, ":::::::::B::*:*W"),
	(0,     0,     1,     'W',     4,     0, ":::::::::B::*:*W"),
	(0,     0,     1,     'W',     0,     0, "::::W::::B::*:*W"),
	(0,     0,     1,     'W',     15,     0, "W:::W::::B::*:*W"),
	(0,     0,     1,     '*',     8,     0, "W:::W::::B::*:*W"),
	(0,     0,     1,     'W',     4,     0, "W:::W:::*B::*:*W"),
	(0,     1,     0,     'B',     0,     0, "W:::W:::*B::*:*W"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, ":*::::::::::::::"),
	(0,     1,     1,     '*',     5,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     9,     0, ":::::*::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::::*::::::*:::"),
	(0,     0,     0,     '*',     8,     0, ":::::*::::::*:::"),
	(0,     0,     0,     'W',     15,     0, ":::::*::::::*:::"),
	(0,     1,     0,     ':',     8,     0, ":::::*::::::*:::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     0,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     3,     0, "::::::W:::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::W::W:::::::::"),
	(0,     0,     1,     'B',     1,     0, ":::W::W:::::::::"),
	(0,     0,     1,     '*',     12,     0, ":B:W::W:::::::::"),
	(0,     0,     0,     'B',     0,     0, ":B:W::W:::::*:::"),
	(0,     0,     0,     'W',     3,     0, ":B:W::W:::::*:::"),
	(0,     0,     1,     'W',     11,     0, ":B:W::W:::::*:::"),
	(0,     0,     1,     '*',     11,     0, ":B:W::W::::W*:::"),
	(0,     0,     0,     ':',     7,     0, ":B:W::W::::B*:::"),
	(0,     0,     1,     'B',     0,     0, ":B:W::W::::B*:::"),
	(0,     0,     0,     'W',     6,     0, "BB:W::W::::B*:::"),
	(0,     0,     1,     ':',     10,     0, "BB:W::W::::B*:::"),
	(0,     0,     0,     '*',     15,     0, "BB:W::W::::B*:::"),
	(0,     0,     1,     '*',     3,     0, "BB:W::W::::B*:::"),
	(0,     1,     0,     ':',     13,     0, "BB:B::W::::B*:::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     10,     0, ":::B::::::::::::"),
	(0,     0,     0,     ':',     13,     0, ":::B::::::::::::"),
	(0,     0,     0,     'B',     5,     0, ":::B::::::::::::"),
	(0,     0,     1,     '*',     15,     0, ":::B::::::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::B:::::::::::*"),
	(0,     0,     0,     'B',     12,     0, ":::B:::::::::::*"),
	(0,     0,     0,     'B',     4,     0, ":::B:::::::::::*"),
	(0,     0,     1,     'B',     0,     0, ":::B:::::::::::*"),
	(0,     0,     1,     ':',     9,     0, "B::B:::::::::::*"),
	(0,     0,     1,     ':',     4,     0, "B::B:::::::::::*"),
	(0,     0,     1,     ':',     11,     0, "B::B:::::::::::*"),
	(0,     1,     0,     '*',     3,     0, "B::B:::::::::::*"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     0, "::::::W:::::::::"),
	(0,     1,     1,     ':',     0,     0, "::::::W:::::::::"),
	(0,     0,     1,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     0, ":::::::::::::*::"),
	(0,     0,     0,     ':',     15,     0, ":::::::::::::*::"),
	(0,     0,     1,     'B',     5,     0, ":::::::::::::*::"),
	(0,     0,     0,     'B',     2,     0, ":::::B:::::::*::"),
	(0,     0,     1,     '*',     11,     0, ":::::B:::::::*::"),
	(0,     0,     0,     'B',     12,     0, ":::::B:::::*:*::"),
	(0,     1,     1,     'W',     9,     0, ":::::B:::::*:*::"),
	(0,     0,     1,     ':',     12,     0, ":::::::::W::::::"),
	(0,     0,     0,     '*',     3,     0, ":::::::::W::::::"),
	(0,     1,     1,     ':',     12,     0, ":::::::::W::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     0, "::::::*:::::::::"),
	(0,     0,     0,     'B',     0,     0, "::::::B:::::::::"),
	(0,     0,     1,     '*',     10,     0, "::::::B:::::::::"),
	(0,     0,     0,     ':',     7,     0, "::::::B:::*:::::"),
	(0,     1,     0,     'B',     6,     0, "::::::B:::*:::::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::*::::::"),
	(0,     0,     1,     'B',     2,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     7,     0, "::B::::::*::::::"),
	(0,     0,     0,     ':',     1,     0, "::B::::::*::::::"),
	(0,     0,     1,     'W',     13,     0, "::B::::::*::::::"),
	(0,     1,     1,     'B',     5,     0, "::B::::::*:::W::"),
	(0,     0,     0,     'B',     6,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     11,     0, ":::::B::::::::::"),
	(0,     0,     0,     'W',     0,     0, ":::::B:::::*::::"),
	(0,     0,     1,     '*',     14,     0, ":::::B:::::*::::"),
	(0,     1,     1,     '*',     14,     0, ":::::B:::::*::*:"),
	(0,     0,     1,     '*',     6,     0, "::::::::::::::*:"),
	(0,     0,     1,     'W',     5,     0, "::::::*:::::::*:"),
	(0,     1,     1,     'B',     7,     0, ":::::W*:::::::*:"),
	(0,     0,     1,     ':',     14,     0, ":::::::B::::::::"),
	(0,     0,     1,     'W',     3,     0, ":::::::B::::::::"),
	(0,     0,     1,     '*',     3,     0, ":::W:::B::::::::"),
	(0,     0,     1,     '*',     9,     0, ":::B:::B::::::::"),
	(0,     0,     0,     'B',     5,     0, ":::B:::B:*::::::"),
	(0,     0,     1,     'W',     13,     0, ":::B:::B:*::::::"),
	(0,     0,     1,     '*',     12,     0, ":::B:::B:*:::W::"),
	(0,     0,     0,     'B',     15,     0, ":::B:::B:*::*W::"),
	(0,     0,     1,     'W',     11,     0, ":::B:::B:*::*W::"),
	(0,     0,     0,     'W',     9,     0, ":::B:::B:*:W*W::"),
	(0,     0,     1,     'W',     15,     0, ":::B:::B:*:W*W::"),
	(0,     0,     0,     ':',     3,     0, ":::B:::B:*:W*W:W"),
	(0,     0,     1,     'W',     12,     0, ":::B:::B:*:W*W:W"),
	(0,     1,     0,     'W',     15,     0, ":::B:::B:*:WWW:W"),
	(0,     1,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     0, ":W::::::::::::::"),
	(0,     0,     1,     'W',     2,     0, ":W:::::::::::B::"),
	(0,     0,     0,     '*',     4,     0, ":WW::::::::::B::"),
	(0,     0,     1,     ':',     0,     0, ":WW::::::::::B::"),
	(1,     0,     1,     ':',     15,     0, ":WW::::::::::B::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     0, "::::::::::B:::::"),
	(0,     0,     0,     'W',     3,     0, "::::::::::B:::::"),
	(0,     0,     1,     '*',     6,     0, "::::::::::B:::::"),
	(0,     1,     1,     ':',     2,     0, "::::::*:::B:::::"),
	(0,     0,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::W:::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::*:W:::::::::::"),
	(0,     0,     1,     'W',     15,     0, "::*:W:::::::::W:"),
	(0,     1,     1,     'B',     7,     0, "::*:W:::::::::WW"),
	(0,     0,     1,     'W',     5,     0, ":::::::B::::::::"),
	(0,     0,     0,     'W',     5,     0, ":::::W:B::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::::W:B::::::::"),
	(0,     0,     1,     'B',     1,     0, ":::::W:B::::::::"),
	(0,     0,     1,     'W',     4,     0, ":B:::W:B::::::::"),
	(0,     0,     1,     '*',     0,     0, ":B::WW:B::::::::"),
	(0,     0,     0,     'B',     2,     0, "*B::WW:B::::::::"),
	(0,     0,     1,     '*',     2,     0, "*B::WW:B::::::::"),
	(0,     0,     1,     ':',     2,     0, "*B*:WW:B::::::::"),
	(0,     0,     1,     'B',     14,     0, "*B*:WW:B::::::::"),
	(0,     0,     0,     ':',     8,     0, "*B*:WW:B::::::B:"),
	(0,     0,     1,     ':',     8,     0, "*B*:WW:B::::::B:"),
	(0,     1,     1,     ':',     12,     0, "*B*:WW:B::::::B:"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::::::*:::::"),
	(0,     0,     0,     'B',     13,     0, "::::::::::*:::::"),
	(0,     0,     0,     ':',     15,     0, "::::::::::*:::::"),
	(0,     0,     0,     'W',     0,     0, "::::::::::*:::::"),
	(0,     0,     1,     'W',     2,     0, "::::::::::*:::::"),
	(0,     0,     1,     'W',     7,     0, "::W:::::::*:::::"),
	(0,     0,     0,     ':',     0,     0, "::W::::W::*:::::"),
	(0,     0,     0,     ':',     10,     0, "::W::::W::*:::::"),
	(0,     0,     1,     'W',     9,     0, "::W::::W::*:::::"),
	(0,     0,     1,     'B',     7,     0, "::W::::W:W*:::::"),
	(0,     1,     0,     ':',     8,     0, "::W::::B:W*:::::"),
	(0,     1,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::::::::::*::"),
	(0,     0,     0,     '*',     1,     0, ":::::::::::::*::"),
	(0,     0,     1,     'B',     9,     0, ":::::::::::::*::"),
	(0,     0,     0,     '*',     8,     0, ":::::::::B:::*::"),
	(0,     0,     0,     ':',     7,     0, ":::::::::B:::*::"),
	(0,     0,     0,     'W',     4,     0, ":::::::::B:::*::"),
	(0,     0,     1,     '*',     4,     0, ":::::::::B:::*::"),
	(0,     0,     0,     'B',     7,     0, "::::*::::B:::*::"),
	(0,     0,     0,     'W',     6,     0, "::::*::::B:::*::"),
	(0,     0,     0,     '*',     0,     0, "::::*::::B:::*::"),
	(0,     0,     1,     'W',     4,     0, "::::*::::B:::*::"),
	(0,     0,     1,     ':',     0,     0, "::::W::::B:::*::"),
	(0,     1,     1,     'W',     15,     0, "::::W::::B:::*::"),
	(0,     0,     0,     ':',     14,     0, ":::::::::::::::W"),
	(0,     0,     1,     '*',     14,     0, ":::::::::::::::W"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::::*W"),
	(0,     0,     0,     '*',     2,     0, "::::::::::::::*W"),
	(0,     1,     1,     ':',     8,     0, "::::::::::::::*W"),
	(1,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, "::::::::::W:::::"),
	(0,     0,     1,     'B',     2,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     12,     0, "::B:::::::W:::::"),
	(0,     1,     1,     '*',     13,     0, "::B:::::::W:::::"),
	(0,     0,     0,     'B',     5,     0, ":::::::::::::*::"),
	(0,     0,     0,     'B',     9,     0, ":::::::::::::*::"),
	(0,     0,     1,     'B',     0,     0, ":::::::::::::*::"),
	(0,     0,     0,     ':',     11,     0, "B::::::::::::*::"),
	(0,     0,     0,     ':',     9,     0, "B::::::::::::*::"),
	(0,     0,     0,     ':',     15,     0, "B::::::::::::*::"),
	(0,     0,     0,     '*',     4,     0, "B::::::::::::*::"),
	(0,     0,     1,     'W',     7,     0, "B::::::::::::*::"),
	(0,     0,     0,     '*',     8,     0, "B::::::W:::::*::"),
	(0,     0,     1,     'B',     5,     0, "B::::::W:::::*::"),
	(0,     0,     0,     '*',     8,     0, "B::::B:W:::::*::"),
	(0,     0,     0,     'B',     7,     0, "B::::B:W:::::*::"),
	(0,     0,     0,     '*',     12,     0, "B::::B:W:::::*::"),
	(0,     0,     0,     'B',     13,     0, "B::::B:W:::::*::"),
	(0,     0,     0,     'W',     15,     0, "B::::B:W:::::*::"),
	(0,     0,     1,     'B',     11,     0, "B::::B:W:::::*::"),
	(0,     0,     1,     'B',     4,     0, "B::::B:W:::B:*::"),
	(0,     0,     0,     '*',     4,     0, "B:::BB:W:::B:*::"),
	(0,     0,     1,     '*',     6,     0, "B:::BB:W:::B:*::"),
	(0,     0,     1,     ':',     7,     0, "B:::BB*W:::B:*::"),
	(0,     0,     0,     '*',     1,     0, "B:::BB*W:::B:*::"),
	(0,     0,     1,     '*',     4,     0, "B:::BB*W:::B:*::"),
	(0,     0,     0,     '*',     2,     0, "B:::WB*W:::B:*::"),
	(0,     0,     1,     ':',     1,     0, "B:::WB*W:::B:*::"),
	(0,     0,     1,     ':',     12,     0, "B:::WB*W:::B:*::"),
	(0,     0,     1,     '*',     14,     0, "B:::WB*W:::B:*::"),
	(0,     0,     1,     ':',     7,     0, "B:::WB*W:::B:**:"),
	(0,     0,     0,     'B',     15,     0, "B:::WB*W:::B:**:"),
	(0,     0,     1,     'W',     3,     0, "B:::WB*W:::B:**:"),
	(0,     0,     0,     '*',     3,     0, "B::WWB*W:::B:**:"),
	(0,     0,     0,     '*',     3,     0, "B::WWB*W:::B:**:"),
	(0,     0,     0,     ':',     15,     0, "B::WWB*W:::B:**:"),
	(0,     0,     0,     'W',     13,     0, "B::WWB*W:::B:**:"),
	(0,     1,     0,     'W',     2,     0, "B::WWB*W:::B:**:"),
	(0,     0,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     1,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     13,     0, ":::::::::::B::::"),
	(0,     1,     0,     '*',     10,     0, ":::::::::::B:*::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":W::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":W::::::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":W::::::::::::::"),
	(0,     1,     0,     ':',     12,     0, ":W:::::::::::*::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(1,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(1,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "::*:::::::::::::"),
	(0,     1,     1,     'W',     12,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     0,     0, "::::::::::::W:::"),
	(0,     0,     0,     'W',     4,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     1,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     1,     0, ":*::::::::::W:::"),
	(0,     0,     0,     '*',     13,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     10,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     14,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     12,     0, "::::::::::::W:W:"),
	(0,     0,     0,     '*',     9,     0, "::::::::::::W:W:"),
	(0,     1,     1,     'B',     13,     0, "::::::::::::W:W:"),
	(0,     0,     0,     '*',     1,     0, ":::::::::::::B::"),
	(0,     0,     0,     '*',     7,     0, ":::::::::::::B::"),
	(0,     0,     0,     'B',     3,     0, ":::::::::::::B::"),
	(0,     0,     0,     '*',     1,     0, ":::::::::::::B::"),
	(0,     1,     1,     'B',     15,     0, ":::::::::::::B::"),
	(0,     0,     1,     '*',     10,     0, ":::::::::::::::B"),
	(0,     0,     0,     'B',     13,     0, "::::::::::*::::B"),
	(0,     0,     1,     'B',     3,     0, "::::::::::*::::B"),
	(0,     0,     1,     ':',     7,     0, ":::B::::::*::::B"),
	(0,     0,     1,     ':',     12,     0, ":::B::::::*::::B"),
	(0,     0,     0,     'B',     4,     0, ":::B::::::*::::B"),
	(0,     0,     1,     'B',     13,     0, ":::B::::::*::::B"),
	(0,     0,     0,     'W',     5,     0, ":::B::::::*::B:B"),
	(0,     0,     0,     '*',     14,     0, ":::B::::::*::B:B"),
	(0,     0,     0,     ':',     6,     0, ":::B::::::*::B:B"),
	(0,     0,     1,     'B',     14,     0, ":::B::::::*::B:B"),
	(0,     1,     0,     'B',     7,     0, ":::B::::::*::BBB"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     0, ":::::::::::B::::"),
	(0,     0,     1,     ':',     1,     0, "::::*::::::B::::"),
	(0,     0,     0,     'W',     8,     0, "::::*::::::B::::"),
	(0,     0,     1,     'W',     12,     0, "::::*::::::B::::"),
	(0,     1,     1,     '*',     12,     0, "::::*::::::BW:::"),
	(0,     0,     0,     '*',     0,     0, "::::::::::::*:::"),
	(0,     0,     1,     '*',     10,     0, "::::::::::::*:::"),
	(0,     0,     0,     'W',     12,     0, "::::::::::*:*:::"),
	(0,     0,     1,     'B',     10,     0, "::::::::::*:*:::"),
	(0,     0,     1,     '*',     4,     0, "::::::::::B:*:::"),
	(0,     0,     0,     '*',     6,     0, "::::*:::::B:*:::"),
	(0,     0,     1,     'W',     9,     0, "::::*:::::B:*:::"),
	(0,     1,     1,     'W',     10,     0, "::::*::::WB:*:::"),
	(0,     0,     1,     'W',     12,     0, "::::::::::W:::::"),
	(0,     0,     1,     ':',     10,     0, "::::::::::W:W:::"),
	(0,     0,     0,     ':',     2,     0, "::::::::::W:W:::"),
	(0,     0,     0,     '*',     3,     0, "::::::::::W:W:::"),
	(0,     0,     0,     'W',     14,     0, "::::::::::W:W:::"),
	(0,     0,     0,     ':',     12,     0, "::::::::::W:W:::"),
	(0,     1,     0,     '*',     9,     0, "::::::::::W:W:::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     0, ":*::::::::::::::"),
	(0,     1,     0,     'B',     2,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "W:::::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "W:::::::::::::::"),
	(0,     0,     0,     'B',     13,     0, "W:::::::::::::::"),
	(0,     0,     0,     'B',     9,     0, "W:::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "W:::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "W:::W:::::::::::"),
	(0,     0,     0,     ':',     6,     0, "W:::W:::::::::::"),
	(0,     0,     0,     '*',     4,     0, "W:::W:::::::::::"),
	(0,     0,     0,     ':',     8,     0, "W:::W:::::::::::"),
	(0,     0,     0,     '*',     11,     0, "W:::W:::::::::::"),
	(0,     0,     0,     ':',     15,     0, "W:::W:::::::::::"),
	(0,     0,     1,     'B',     13,     0, "W:::W:::::::::::"),
	(0,     0,     1,     ':',     5,     0, "W:::W::::::::B::"),
	(0,     0,     1,     'B',     5,     0, "W:::W::::::::B::"),
	(0,     0,     0,     'W',     13,     0, "W:::WB:::::::B::"),
	(0,     0,     1,     'W',     1,     0, "W:::WB:::::::B::"),
	(0,     0,     1,     ':',     10,     0, "WW::WB:::::::B::"),
	(0,     1,     0,     'B',     4,     0, "WW::WB:::::::B::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     13,     0, "::::::::::::::B:"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     14,     0, ":::::B:::::W::::"),
	(0,     0,     0,     '*',     8,     0, ":::::B:::::W::B:"),
	(0,     0,     1,     ':',     3,     0, ":::::B:::::W::B:"),
	(0,     0,     1,     'W',     6,     0, ":::::B:::::W::B:"),
	(0,     1,     1,     '*',     3,     0, ":::::BW::::W::B:"),
	(0,     0,     1,     ':',     4,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     15,     0, ":::*::::::::::::"),
	(0,     0,     1,     'W',     10,     0, ":::*::::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::*::::::W:::::"),
	(0,     0,     0,     ':',     4,     0, ":::*::::::W:::W:"),
	(0,     0,     0,     'W',     11,     0, ":::*::::::W:::W:"),
	(0,     0,     1,     '*',     8,     0, ":::*::::::W:::W:"),
	(0,     0,     0,     '*',     15,     0, ":::*::::*:W:::W:"),
	(0,     0,     0,     '*',     10,     0, ":::*::::*:W:::W:"),
	(0,     0,     0,     'W',     4,     0, ":::*::::*:W:::W:"),
	(0,     0,     1,     '*',     0,     0, ":::*::::*:W:::W:"),
	(0,     0,     0,     '*',     3,     0, "*::*::::*:W:::W:"),
	(0,     0,     0,     '*',     5,     0, "*::*::::*:W:::W:"),
	(0,     0,     1,     'W',     10,     0, "*::*::::*:W:::W:"),
	(0,     0,     1,     'W',     5,     0, "*::*::::*:W:::W:"),
	(0,     0,     1,     'W',     0,     0, "*::*:W::*:W:::W:"),
	(0,     0,     1,     ':',     5,     0, "W::*:W::*:W:::W:"),
	(0,     0,     0,     '*',     5,     0, "W::*:W::*:W:::W:"),
	(0,     0,     0,     ':',     12,     0, "W::*:W::*:W:::W:"),
	(0,     0,     1,     'B',     8,     0, "W::*:W::*:W:::W:"),
	(0,     0,     1,     '*',     10,     0, "W::*:W::B:W:::W:"),
	(0,     0,     1,     'W',     13,     0, "W::*:W::B:B:::W:"),
	(0,     0,     1,     ':',     13,     0, "W::*:W::B:B::WW:"),
	(0,     0,     1,     'W',     15,     0, "W::*:W::B:B::WW:"),
	(0,     0,     1,     ':',     13,     0, "W::*:W::B:B::WWW"),
	(0,     0,     1,     '*',     4,     0, "W::*:W::B:B::WWW"),
	(0,     0,     0,     ':',     12,     0, "W::**W::B:B::WWW"),
	(0,     0,     0,     'W',     10,     0, "W::**W::B:B::WWW"),
	(0,     0,     1,     '*',     0,     0, "W::**W::B:B::WWW"),
	(0,     0,     1,     ':',     10,     0, "B::**W::B:B::WWW"),
	(0,     0,     0,     ':',     14,     0, "B::**W::B:B::WWW"),
	(0,     0,     0,     'W',     9,     0, "B::**W::B:B::WWW"),
	(0,     0,     1,     ':',     8,     0, "B::**W::B:B::WWW"),
	(0,     0,     0,     '*',     15,     0, "B::**W::B:B::WWW"),
	(0,     0,     0,     'B',     14,     0, "B::**W::B:B::WWW"),
	(0,     0,     1,     'W',     8,     0, "B::**W::B:B::WWW"),
	(0,     1,     1,     '*',     13,     0, "B::**W::W:B::WWW"),
	(0,     0,     0,     ':',     0,     0, ":::::::::::::*::"),
	(0,     1,     1,     ':',     0,     0, ":::::::::::::*::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::::*::::::::"),
	(0,     0,     1,     'B',     14,     0, ":::::::*::::::::"),
	(0,     1,     1,     '*',     13,     0, ":::::::*::::::B:"),
	(0,     0,     0,     '*',     8,     0, ":::::::::::::*::"),
	(0,     0,     0,     'W',     4,     0, ":::::::::::::*::"),
	(0,     0,     0,     'W',     4,     0, ":::::::::::::*::"),
	(0,     1,     0,     ':',     4,     0, ":::::::::::::*::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     3,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::*:::::::::::::"),
	(0,     1,     0,     'B',     10,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     0, "W:::::::::::::::"),
	(0,     0,     1,     ':',     3,     0, "W::::::*::::::::"),
	(0,     0,     0,     ':',     2,     0, "W::::::*::::::::"),
	(0,     0,     0,     'B',     8,     0, "W::::::*::::::::"),
	(0,     0,     0,     'W',     10,     0, "W::::::*::::::::"),
	(0,     0,     1,     'B',     9,     0, "W::::::*::::::::"),
	(0,     0,     0,     ':',     10,     0, "W::::::*:B::::::"),
	(0,     0,     1,     '*',     1,     0, "W::::::*:B::::::"),
	(0,     0,     0,     'B',     12,     0, "W*:::::*:B::::::"),
	(0,     0,     0,     'W',     3,     0, "W*:::::*:B::::::"),
	(0,     0,     0,     '*',     7,     0, "W*:::::*:B::::::"),
	(0,     0,     0,     '*',     7,     0, "W*:::::*:B::::::"),
	(0,     0,     1,     'B',     3,     0, "W*:::::*:B::::::"),
	(0,     0,     0,     'B',     13,     0, "W*:B:::*:B::::::"),
	(0,     0,     0,     'W',     11,     0, "W*:B:::*:B::::::"),
	(0,     0,     1,     'B',     7,     0, "W*:B:::*:B::::::"),
	(0,     1,     0,     '*',     2,     0, "W*:B:::B:B::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     14,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     12,     0, "::::::W:::::::W:"),
	(1,     0,     0,     'W',     11,     0, "::::::W:::::::W:"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     0, "::::*:::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::*::::::::B::"),
	(0,     0,     0,     'B',     2,     0, "::::*::::::::B::"),
	(0,     0,     0,     'W',     12,     0, "::::*::::::::B::"),
	(0,     0,     0,     'B',     7,     0, "::::*::::::::B::"),
	(0,     1,     0,     '*',     3,     0, "::::*::::::::B::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     0, "*:::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, "*:::B:::::::::::"),
	(0,     0,     0,     'W',     8,     0, "*:::B:::::::::::"),
	(0,     0,     1,     ':',     8,     0, "*:::B:::::::::::"),
	(0,     0,     0,     '*',     1,     0, "*:::B:::::::::::"),
	(0,     0,     1,     'W',     6,     0, "*:::B:::::::::::"),
	(0,     0,     1,     'B',     12,     0, "*:::B:W:::::::::"),
	(0,     0,     1,     'B',     12,     0, "*:::B:W:::::B:::"),
	(0,     0,     0,     'W',     13,     0, "*:::B:W:::::B:::"),
	(0,     0,     0,     ':',     10,     0, "*:::B:W:::::B:::"),
	(0,     0,     0,     'B',     1,     0, "*:::B:W:::::B:::"),
	(0,     0,     1,     '*',     15,     0, "*:::B:W:::::B:::"),
	(0,     0,     0,     'W',     11,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     'W',     6,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     '*',     14,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     '*',     10,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     'W',     9,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     ':',     5,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     '*',     5,     0, "*:::B:W:::::B::*"),
	(0,     0,     0,     '*',     10,     0, "*:::B:W:::::B::*"),
	(0,     0,     1,     '*',     9,     0, "*:::B:W:::::B::*"),
	(0,     0,     1,     '*',     8,     0, "*:::B:W::*::B::*"),
	(0,     0,     0,     ':',     3,     0, "*:::B:W:**::B::*"),
	(0,     0,     1,     'W',     6,     0, "*:::B:W:**::B::*"),
	(0,     0,     0,     '*',     2,     0, "*:::B:W:**::B::*"),
	(0,     0,     0,     'W',     0,     0, "*:::B:W:**::B::*"),
	(0,     0,     1,     ':',     6,     0, "*:::B:W:**::B::*"),
	(0,     0,     1,     'B',     15,     0, "*:::B:W:**::B::*"),
	(0,     1,     1,     '*',     1,     0, "*:::B:W:**::B::B"),
	(0,     0,     0,     'B',     5,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     15,     0, ":*::::::::::::::"),
	(1,     1,     1,     'W',     3,     0, ":*:::::::::::::B"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(1,     0,     0,     '*',     6,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     0, ":::::::::::::::B"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     10,     0, ":::::::::::::::B"),
	(0,     0,     1,     '*',     14,     0, ":::::::::::::::B"),
	(0,     0,     1,     'B',     2,     0, "::::::::::::::*B"),
	(0,     0,     1,     '*',     7,     0, "::B:::::::::::*B"),
	(0,     0,     0,     ':',     3,     0, "::B::::*::::::*B"),
	(0,     0,     1,     '*',     8,     0, "::B::::*::::::*B"),
	(0,     0,     0,     '*',     1,     0, "::B::::**:::::*B"),
	(0,     0,     0,     'W',     8,     0, "::B::::**:::::*B"),
	(0,     0,     0,     ':',     5,     0, "::B::::**:::::*B"),
	(0,     0,     1,     '*',     2,     0, "::B::::**:::::*B"),
	(0,     0,     0,     '*',     10,     0, "::W::::**:::::*B"),
	(0,     0,     0,     '*',     2,     0, "::W::::**:::::*B"),
	(0,     0,     0,     '*',     10,     0, "::W::::**:::::*B"),
	(0,     0,     1,     'W',     8,     0, "::W::::**:::::*B"),
	(0,     0,     1,     ':',     11,     0, "::W::::*W:::::*B"),
	(0,     0,     1,     'B',     15,     0, "::W::::*W:::::*B"),
	(0,     1,     1,     '*',     15,     0, "::W::::*W:::::*B"),
	(0,     0,     0,     'W',     5,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     1,     0, ":::::::::::::::*"),
	(0,     0,     1,     ':',     10,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     10,     0, ":::::::::::::::*"),
	(0,     0,     0,     'W',     12,     0, ":::::::::::::::*"),
	(0,     0,     0,     'W',     13,     0, ":::::::::::::::*"),
	(0,     0,     1,     'B',     4,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     3,     0, "::::B::::::::::*"),
	(0,     0,     1,     ':',     10,     0, "::::B::::::::::*"),
	(0,     0,     0,     '*',     2,     0, "::::B::::::::::*"),
	(0,     0,     0,     ':',     4,     0, "::::B::::::::::*"),
	(0,     0,     1,     ':',     10,     0, "::::B::::::::::*"),
	(0,     0,     0,     'W',     3,     0, "::::B::::::::::*"),
	(0,     0,     1,     '*',     2,     0, "::::B::::::::::*"),
	(0,     0,     1,     '*',     14,     0, "::*:B::::::::::*"),
	(0,     1,     0,     'B',     15,     0, "::*:B:::::::::**"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     0, "::::::::::*:::::"),
	(0,     0,     1,     'B',     10,     0, "::::::::::*:::::"),
	(0,     0,     0,     ':',     10,     0, "::::::::::B:::::"),
	(0,     0,     1,     '*',     6,     0, "::::::::::B:::::"),
	(0,     0,     0,     'B',     14,     0, "::::::*:::B:::::"),
	(0,     0,     0,     'W',     9,     0, "::::::*:::B:::::"),
	(0,     0,     0,     'B',     2,     0, "::::::*:::B:::::"),
	(0,     0,     1,     'W',     13,     0, "::::::*:::B:::::"),
	(0,     0,     0,     ':',     3,     0, "::::::*:::B::W::"),
	(0,     0,     0,     ':',     13,     0, "::::::*:::B::W::"),
	(0,     0,     0,     'B',     11,     0, "::::::*:::B::W::"),
	(0,     0,     0,     ':',     11,     0, "::::::*:::B::W::"),
	(0,     0,     0,     ':',     11,     0, "::::::*:::B::W::"),
	(0,     0,     0,     ':',     6,     0, "::::::*:::B::W::"),
	(0,     0,     1,     ':',     7,     0, "::::::*:::B::W::"),
	(0,     0,     1,     'W',     2,     0, "::::::*:::B::W::"),
	(0,     0,     0,     'B',     5,     0, "::W:::*:::B::W::"),
	(0,     0,     0,     'B',     8,     0, "::W:::*:::B::W::"),
	(0,     0,     1,     ':',     7,     0, "::W:::*:::B::W::"),
	(0,     0,     1,     ':',     3,     0, "::W:::*:::B::W::"),
	(0,     0,     0,     ':',     12,     0, "::W:::*:::B::W::"),
	(0,     0,     1,     ':',     12,     0, "::W:::*:::B::W::"),
	(0,     0,     0,     'W',     0,     0, "::W:::*:::B::W::"),
	(0,     0,     0,     '*',     9,     0, "::W:::*:::B::W::"),
	(0,     0,     1,     'B',     3,     0, "::W:::*:::B::W::"),
	(0,     0,     1,     'B',     1,     0, "::WB::*:::B::W::"),
	(0,     0,     1,     'B',     10,     0, ":BWB::*:::B::W::"),
	(0,     0,     0,     'W',     14,     0, ":BWB::*:::B::W::"),
	(0,     0,     0,     '*',     12,     0, ":BWB::*:::B::W::"),
	(0,     0,     1,     ':',     8,     0, ":BWB::*:::B::W::"),
	(0,     1,     1,     ':',     0,     0, ":BWB::*:::B::W::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     0, "::::::::::::*:::"),
	(0,     0,     1,     ':',     8,     0, "::::::::::::*:::"),
	(0,     0,     0,     'W',     10,     0, "::::::::::::*:::"),
	(0,     0,     0,     'W',     15,     0, "::::::::::::*:::"),
	(0,     1,     0,     ':',     7,     0, "::::::::::::*:::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     0, "::::::::::::B:::"),
	(0,     0,     1,     '*',     5,     0, "::::::::::::B:::"),
	(0,     0,     0,     'W',     10,     0, ":::::*::::::B:::"),
	(0,     0,     1,     ':',     0,     0, ":::::*::::::B:::"),
	(0,     0,     1,     ':',     15,     0, ":::::*::::::B:::"),
	(0,     0,     1,     ':',     8,     0, ":::::*::::::B:::"),
	(0,     0,     0,     'B',     8,     0, ":::::*::::::B:::"),
	(0,     0,     1,     'W',     0,     0, ":::::*::::::B:::"),
	(0,     0,     1,     ':',     12,     0, "W::::*::::::B:::"),
	(0,     1,     1,     ':',     12,     0, "W::::*::::::B:::"),
	(0,     1,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, "::::*:::::::::::"),
	(0,     1,     1,     'W',     4,     0, "::::*::::::B::::"),
	(0,     0,     0,     ':',     9,     0, "::::W:::::::::::"),
	(0,     0,     0,     ':',     12,     0, "::::W:::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::::W:::::::::::"),
	(0,     0,     0,     'W',     15,     0, "::::W:::::::::::"),
	(0,     1,     0,     'B',     8,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     0, "B:::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, "B:::::::::::::::"),
	(0,     0,     0,     'B',     9,     0, "B::::::::::W::::"),
	(0,     0,     0,     ':',     14,     0, "B::::::::::W::::"),
	(0,     1,     0,     ':',     12,     0, "B::::::::::W::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     11,     0, ":::::::::::W::::"),
	(0,     0,     0,     ':',     6,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     13,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     0,     0, ":::::::::::B::::"),
	(0,     0,     1,     'W',     15,     0, "*::::::::::B::::"),
	(0,     1,     0,     'W',     4,     0, "*::::::::::B:::W"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     0,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, "::::::::::::B:::"),
	(0,     0,     0,     ':',     13,     0, "::::::::::::B:::"),
	(0,     0,     0,     ':',     1,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     3,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     14,     0, ":::W::::::::B:::"),
	(0,     0,     1,     '*',     10,     0, ":::W::::::::B:W:"),
	(0,     0,     0,     'W',     14,     0, ":::W::::::*:B:W:"),
	(0,     0,     1,     ':',     2,     0, ":::W::::::*:B:W:"),
	(0,     1,     0,     ':',     10,     0, ":::W::::::*:B:W:"),
	(0,     1,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, "B:::::::::::::::"),
	(0,     0,     0,     'B',     11,     0, "B:::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, "B:::::::::::::::"),
	(0,     1,     0,     'W',     4,     0, "B::::::::::B::::"),
	(0,     1,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     4,     0, ":::::::B:::W::::"),
	(0,     1,     0,     ':',     8,     0, ":::::::B:::W::::"),
	(0,     0,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     3,     0, "::::W:::::::::::"),
	(0,     0,     0,     'B',     12,     0, ":::WW:::::::::::"),
	(0,     0,     0,     'W',     13,     0, ":::WW:::::::::::"),
	(0,     0,     0,     'B',     8,     0, ":::WW:::::::::::"),
	(1,     0,     1,     '*',     3,     0, ":::WW:::::::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, "::::::*:::::::::"),
	(0,     0,     0,     'W',     3,     0, "::::::*:::::::::"),
	(0,     0,     0,     'B',     1,     0, "::::::*:::::::::"),
	(0,     0,     0,     ':',     8,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     0,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     14,     0, "W:::::*:::::::::"),
	(0,     0,     1,     ':',     2,     0, "W:::::*:::::::::"),
	(0,     0,     1,     ':',     11,     0, "W:::::*:::::::::"),
	(1,     0,     1,     '*',     15,     0, "W:::::*:::::::::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     0, "::::::::B:::::::"),
	(0,     0,     0,     'B',     2,     0, "::::::::B:::::::"),
	(0,     1,     0,     '*',     5,     0, "::::::::B:::::::"),
	(0,     0,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     12,     0, "::::::::::B:::::"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     0, "::::::::::::::B:"),
	(0,     0,     0,     'W',     11,     0, "::::::::::::::B:"),
	(0,     0,     1,     'B',     3,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     11,     0, ":::B::::::::::B:"),
	(0,     0,     0,     ':',     9,     0, ":::B::::::::::B:"),
	(0,     1,     0,     'W',     2,     0, ":::B::::::::::B:"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":*::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     0,     0, "**::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, "**::::::::::::::"),
	(0,     0,     0,     '*',     6,     0, "**::::::::::::::"),
	(0,     0,     1,     'W',     7,     0, "**::::::::::::::"),
	(0,     0,     1,     'W',     5,     0, "**:::::W::::::::"),
	(0,     0,     0,     'W',     12,     0, "**:::W:W::::::::"),
	(0,     0,     0,     'W',     2,     0, "**:::W:W::::::::"),
	(0,     0,     0,     'B',     10,     0, "**:::W:W::::::::"),
	(0,     0,     0,     '*',     12,     0, "**:::W:W::::::::"),
	(0,     0,     1,     'B',     5,     0, "**:::W:W::::::::"),
	(0,     0,     1,     ':',     2,     0, "**:::B:W::::::::"),
	(0,     0,     1,     'W',     6,     0, "**:::B:W::::::::"),
	(0,     0,     1,     ':',     1,     0, "**:::BWW::::::::"),
	(0,     0,     1,     'W',     5,     0, "**:::BWW::::::::"),
	(0,     0,     0,     'B',     9,     0, "**:::WWW::::::::"),
	(0,     0,     1,     '*',     1,     0, "**:::WWW::::::::"),
	(0,     0,     0,     '*',     8,     0, "*::::WWW::::::::"),
	(0,     0,     1,     'B',     4,     0, "*::::WWW::::::::"),
	(0,     0,     0,     ':',     0,     0, "*:::BWWW::::::::"),
	(0,     0,     1,     ':',     0,     0, "*:::BWWW::::::::"),
	(0,     0,     1,     'W',     5,     0, "*:::BWWW::::::::"),
	(0,     0,     1,     ':',     15,     0, "*:::BWWW::::::::"),
	(0,     0,     1,     'W',     7,     0, "*:::BWWW::::::::"),
	(0,     0,     1,     'W',     6,     0, "*:::BWWW::::::::"),
	(0,     0,     0,     'W',     8,     0, "*:::BWWW::::::::"),
	(0,     0,     0,     '*',     2,     0, "*:::BWWW::::::::"),
	(0,     0,     0,     '*',     5,     0, "*:::BWWW::::::::"),
	(0,     1,     0,     ':',     13,     0, "*:::BWWW::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     0, "::B:::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "::B:::::::::::::"),
	(0,     0,     1,     ':',     11,     0, "::B:::::::::::::"),
	(0,     0,     1,     ':',     0,     0, "::B:::::::::::::"),
	(0,     0,     0,     '*',     7,     0, "::B:::::::::::::"),
	(0,     1,     1,     ':',     14,     0, "::B:::::::::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     0, ":::::::::::::B::"),
	(0,     1,     1,     'W',     6,     0, ":::::::::*:::B::"),
	(0,     0,     0,     '*',     15,     0, "::::::W:::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     7,     0, "::*:::W:::::::::"),
	(0,     0,     1,     'B',     13,     0, "::*:::W:::::::::"),
	(0,     0,     1,     '*',     4,     0, "::*:::W::::::B::"),
	(0,     0,     0,     'B',     2,     0, "::*:*:W::::::B::"),
	(0,     0,     1,     '*',     15,     0, "::*:*:W::::::B::"),
	(0,     0,     0,     'B',     15,     0, "::*:*:W::::::B:*"),
	(0,     0,     1,     '*',     13,     0, "::*:*:W::::::B:*"),
	(0,     0,     1,     'W',     3,     0, "::*:*:W::::::W:*"),
	(0,     0,     1,     ':',     1,     0, "::*W*:W::::::W:*"),
	(0,     0,     1,     'B',     1,     0, "::*W*:W::::::W:*"),
	(0,     1,     0,     ':',     6,     0, ":B*W*:W::::::W:*"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     0, "*:::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, "*:::::::::::::::"),
	(0,     0,     1,     '*',     6,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     13,     0, "*:::::*:::::::::"),
	(0,     0,     0,     '*',     13,     0, "*:::::*:::::::::"),
	(0,     0,     1,     '*',     15,     0, "*:::::*:::::::::"),
	(0,     0,     1,     '*',     9,     0, "*:::::*::::::::*"),
	(0,     0,     1,     'B',     10,     0, "*:::::*::*:::::*"),
	(0,     0,     1,     'B',     11,     0, "*:::::*::*B::::*"),
	(0,     0,     0,     'B',     12,     0, "*:::::*::*BB:::*"),
	(0,     1,     0,     ':',     11,     0, "*:::::*::*BB:::*"),
	(0,     0,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     2,     0, "::::::::::B:::::"),
	(0,     0,     0,     '*',     8,     0, "::W:::::::B:::::"),
	(0,     0,     0,     'B',     3,     0, "::W:::::::B:::::"),
	(0,     0,     1,     ':',     15,     0, "::W:::::::B:::::"),
	(0,     0,     0,     '*',     6,     0, "::W:::::::B:::::"),
	(0,     0,     0,     ':',     1,     0, "::W:::::::B:::::"),
	(0,     0,     1,     ':',     14,     0, "::W:::::::B:::::"),
	(0,     0,     0,     'B',     9,     0, "::W:::::::B:::::"),
	(0,     0,     0,     'B',     11,     0, "::W:::::::B:::::"),
	(0,     0,     1,     '*',     6,     0, "::W:::::::B:::::"),
	(0,     0,     0,     'W',     12,     0, "::W:::*:::B:::::"),
	(0,     0,     1,     'W',     7,     0, "::W:::*:::B:::::"),
	(0,     0,     0,     'B',     7,     0, "::W:::*W::B:::::"),
	(0,     0,     1,     'W',     5,     0, "::W:::*W::B:::::"),
	(0,     0,     1,     '*',     2,     0, "::W::W*W::B:::::"),
	(0,     0,     0,     'W',     15,     0, "::B::W*W::B:::::"),
	(0,     0,     0,     '*',     7,     0, "::B::W*W::B:::::"),
	(0,     0,     0,     '*',     13,     0, "::B::W*W::B:::::"),
	(0,     0,     0,     '*',     1,     0, "::B::W*W::B:::::"),
	(0,     0,     1,     '*',     3,     0, "::B::W*W::B:::::"),
	(0,     0,     0,     '*',     10,     0, "::B*:W*W::B:::::"),
	(0,     0,     1,     ':',     3,     0, "::B*:W*W::B:::::"),
	(0,     0,     0,     '*',     12,     0, "::B*:W*W::B:::::"),
	(0,     1,     0,     'W',     11,     0, "::B*:W*W::B:::::"),
	(0,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::::::::::::W:::"),
	(0,     0,     0,     'W',     15,     0, "::::::::::::W:::"),
	(0,     0,     0,     'W',     7,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     5,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     5,     0, ":::::*::::::W:::"),
	(0,     0,     1,     'B',     9,     0, ":::::*::::::W:::"),
	(0,     0,     1,     '*',     8,     0, ":::::*:::B::W:::"),
	(0,     0,     1,     '*',     6,     0, ":::::*::*B::W:::"),
	(0,     0,     0,     ':',     8,     0, ":::::**:*B::W:::"),
	(0,     0,     1,     'B',     1,     0, ":::::**:*B::W:::"),
	(0,     0,     1,     'W',     9,     0, ":B:::**:*B::W:::"),
	(0,     0,     0,     'B',     14,     0, ":B:::**:*W::W:::"),
	(0,     0,     0,     '*',     13,     0, ":B:::**:*W::W:::"),
	(0,     0,     0,     'B',     5,     0, ":B:::**:*W::W:::"),
	(0,     0,     0,     'W',     3,     0, ":B:::**:*W::W:::"),
	(0,     0,     1,     'W',     7,     0, ":B:::**:*W::W:::"),
	(0,     0,     1,     ':',     8,     0, ":B:::**W*W::W:::"),
	(0,     0,     0,     '*',     12,     0, ":B:::**W*W::W:::"),
	(0,     0,     1,     '*',     3,     0, ":B:::**W*W::W:::"),
	(0,     0,     0,     ':',     1,     0, ":B:*:**W*W::W:::"),
	(0,     1,     1,     'W',     14,     0, ":B:*:**W*W::W:::"),
	(0,     0,     0,     '*',     5,     0, "::::::::::::::W:"),
	(0,     0,     1,     '*',     10,     0, "::::::::::::::W:"),
	(0,     0,     1,     'W',     12,     0, "::::::::::*:::W:"),
	(1,     0,     0,     'W',     5,     0, "::::::::::*:W:W:"),
	(0,     1,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     10,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     10,     0, "::::::::::*:::::"),
	(0,     0,     0,     ':',     6,     0, "::::::::::*:::::"),
	(0,     1,     0,     ':',     8,     0, "::::::::::*:::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::::::::*:::::::"),
	(0,     0,     1,     ':',     1,     0, "::::::::*:::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::::*:::::::"),
	(0,     1,     0,     ':',     2,     0, "::::::::*:::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     5,     0, "::*::::::*::::::"),
	(0,     0,     1,     '*',     7,     0, "::*::::::*::::::"),
	(0,     0,     0,     'B',     2,     0, "::*::::*:*::::::"),
	(0,     0,     1,     '*',     10,     0, "::*::::*:*::::::"),
	(0,     0,     0,     'B',     12,     0, "::*::::*:**:::::"),
	(0,     0,     1,     '*',     6,     0, "::*::::*:**:::::"),
	(0,     0,     1,     '*',     15,     0, "::*:::**:**:::::"),
	(0,     0,     1,     'B',     6,     0, "::*:::**:**::::*"),
	(0,     0,     0,     ':',     2,     0, "::*:::B*:**::::*"),
	(0,     0,     1,     '*',     6,     0, "::*:::B*:**::::*"),
	(0,     0,     0,     'B',     5,     0, "::*:::W*:**::::*"),
	(0,     0,     1,     '*',     4,     0, "::*:::W*:**::::*"),
	(0,     0,     1,     'B',     13,     0, "::*:*:W*:**::::*"),
	(0,     0,     1,     'W',     14,     0, "::*:*:W*:**::B:*"),
	(0,     0,     1,     'B',     2,     0, "::*:*:W*:**::BW*"),
	(0,     0,     0,     'W',     2,     0, "::B:*:W*:**::BW*"),
	(0,     0,     1,     ':',     10,     0, "::B:*:W*:**::BW*"),
	(0,     0,     1,     ':',     9,     0, "::B:*:W*:**::BW*"),
	(0,     0,     0,     'B',     0,     0, "::B:*:W*:**::BW*"),
	(0,     0,     1,     'B',     15,     0, "::B:*:W*:**::BW*"),
	(1,     0,     0,     'B',     15,     0, "::B:*:W*:**::BWB"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::W:::::"),
	(0,     0,     0,     ':',     9,     0, "::::::::::W:::::"),
	(0,     0,     1,     'W',     5,     0, "::::::::::W:::::"),
	(0,     0,     0,     ':',     11,     0, ":::::W::::W:::::"),
	(0,     0,     0,     'B',     11,     0, ":::::W::::W:::::"),
	(0,     0,     1,     'B',     3,     0, ":::::W::::W:::::"),
	(0,     0,     0,     'B',     2,     0, ":::B:W::::W:::::"),
	(0,     0,     1,     ':',     1,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     'B',     0,     0, ":::B:W::::W:::::"),
	(0,     0,     1,     ':',     12,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     '*',     11,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     ':',     7,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     ':',     6,     0, ":::B:W::::W:::::"),
	(0,     0,     1,     ':',     14,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     'W',     3,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     '*',     15,     0, ":::B:W::::W:::::"),
	(0,     0,     1,     'B',     9,     0, ":::B:W::::W:::::"),
	(0,     0,     0,     'B',     11,     0, ":::B:W:::BW:::::"),
	(0,     0,     1,     '*',     5,     0, ":::B:W:::BW:::::"),
	(0,     1,     1,     ':',     13,     0, ":::B:B:::BW:::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     2,     0, "::::::B:::::::::"),
	(0,     0,     1,     'B',     12,     0, "::W:::::::::::::"),
	(0,     0,     0,     '*',     0,     0, "::W:::::::::B:::"),
	(0,     0,     1,     ':',     0,     0, "::W:::::::::B:::"),
	(0,     0,     1,     'B',     8,     0, "::W:::::::::B:::"),
	(0,     0,     1,     'B',     13,     0, "::W:::::B:::B:::"),
	(0,     0,     1,     'W',     13,     0, "::W:::::B:::BB::"),
	(0,     0,     1,     '*',     12,     0, "::W:::::B:::BW::"),
	(0,     0,     1,     '*',     7,     0, "::W:::::B:::WW::"),
	(0,     0,     0,     'W',     4,     0, "::W::::*B:::WW::"),
	(0,     0,     0,     '*',     15,     0, "::W::::*B:::WW::"),
	(0,     0,     0,     ':',     2,     0, "::W::::*B:::WW::"),
	(0,     0,     0,     '*',     14,     0, "::W::::*B:::WW::"),
	(0,     0,     1,     '*',     3,     0, "::W::::*B:::WW::"),
	(0,     0,     0,     ':',     12,     0, "::W*:::*B:::WW::"),
	(0,     1,     1,     'W',     2,     0, "::W*:::*B:::WW::"),
	(0,     0,     1,     ':',     13,     0, "::W:::::::::::::"),
	(0,     1,     1,     ':',     3,     0, "::W:::::::::::::"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     8,     0, "::::::::::::::B:"),
	(0,     0,     1,     '*',     2,     0, "::::::::::::::B:"),
	(0,     0,     0,     '*',     7,     0, "::*:::::::::::B:"),
	(0,     0,     0,     ':',     15,     0, "::*:::::::::::B:"),
	(0,     1,     1,     'B',     4,     0, "::*:::::::::::B:"),
	(0,     0,     1,     '*',     7,     0, "::::B:::::::::::"),
	(0,     0,     1,     ':',     1,     0, "::::B::*::::::::"),
	(0,     0,     1,     '*',     6,     0, "::::B::*::::::::"),
	(0,     0,     0,     '*',     9,     0, "::::B:**::::::::"),
	(0,     0,     1,     ':',     0,     0, "::::B:**::::::::"),
	(0,     1,     0,     'B',     4,     0, "::::B:**::::::::"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     0, "W:::::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "W:::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, "W:::::::::::::::"),
	(0,     1,     0,     ':',     12,     0, "W::::::::::::::W"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     0,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     9,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, ":*:::::::B::::::"),
	(0,     0,     1,     '*',     5,     0, ":*:::::::B::::::"),
	(0,     1,     1,     '*',     0,     0, ":*:::*:::B::::::"),
	(0,     0,     0,     'B',     12,     0, "*:::::::::::::::"),
	(0,     0,     1,     ':',     14,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, "*:::::::::::::::"),
	(0,     0,     1,     'W',     8,     0, "*:::::::::::::::"),
	(0,     1,     1,     '*',     3,     0, "*:::::::W:::::::"),
	(0,     0,     0,     ':',     0,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::*::::::::::::"),
	(0,     0,     0,     'B',     9,     0, ":::*::::::::::::"),
	(0,     0,     1,     'W',     8,     0, ":::*::::::::::::"),
	(0,     0,     0,     'B',     15,     0, ":::*::::W:::::::"),
	(0,     1,     0,     '*',     4,     0, ":::*::::W:::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::W::::*::::::"),
	(0,     0,     1,     'B',     2,     0, "::::W::::*B:::::"),
	(0,     0,     1,     '*',     10,     0, "::B:W::::*B:::::"),
	(0,     0,     0,     '*',     8,     0, "::B:W::::*W:::::"),
	(0,     0,     1,     'W',     8,     0, "::B:W::::*W:::::"),
	(0,     0,     0,     '*',     4,     0, "::B:W:::W*W:::::"),
	(0,     0,     0,     ':',     10,     0, "::B:W:::W*W:::::"),
	(0,     0,     0,     'W',     15,     0, "::B:W:::W*W:::::"),
	(0,     0,     1,     ':',     0,     0, "::B:W:::W*W:::::"),
	(0,     0,     1,     'B',     10,     0, "::B:W:::W*W:::::"),
	(0,     0,     1,     ':',     4,     0, "::B:W:::W*B:::::"),
	(0,     0,     1,     'W',     12,     0, "::B:W:::W*B:::::"),
	(0,     0,     1,     'W',     2,     0, "::B:W:::W*B:W:::"),
	(0,     0,     1,     ':',     15,     0, "::W:W:::W*B:W:::"),
	(0,     0,     1,     'B',     14,     0, "::W:W:::W*B:W:::"),
	(0,     0,     1,     '*',     12,     0, "::W:W:::W*B:W:B:"),
	(0,     0,     1,     ':',     10,     0, "::W:W:::W*B:B:B:"),
	(0,     0,     1,     'B',     6,     0, "::W:W:::W*B:B:B:"),
	(0,     1,     1,     'B',     5,     0, "::W:W:B:W*B:B:B:"),
	(0,     0,     0,     '*',     14,     0, ":::::B::::::::::"),
	(0,     0,     1,     'W',     8,     0, ":::::B::::::::::"),
	(0,     0,     1,     'W',     10,     0, ":::::B::W:::::::"),
	(0,     1,     0,     'W',     8,     0, ":::::B::W:W:::::"),
	(0,     1,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     0, "::::B:::::::::::"),
	(0,     0,     0,     '*',     15,     0, "::::BW::::::::::"),
	(0,     0,     0,     ':',     1,     0, "::::BW::::::::::"),
	(0,     0,     0,     'W',     2,     0, "::::BW::::::::::"),
	(0,     0,     1,     ':',     4,     0, "::::BW::::::::::"),
	(0,     0,     1,     'W',     12,     0, "::::BW::::::::::"),
	(0,     0,     0,     ':',     14,     0, "::::BW::::::W:::"),
	(0,     1,     1,     ':',     10,     0, "::::BW::::::W:::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     13,     0, "::::::::::::W:::"),
	(0,     1,     0,     'B',     11,     0, "::::::::::::W:::"),
	(0,     0,     1,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":B::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, ":B::::::::::::::"),
	(0,     1,     1,     '*',     12,     0, ":B:::::::W::::::"),
	(0,     1,     0,     'W',     3,     0, "::::::::::::*:::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::*::::::::::"),
	(0,     0,     1,     'B',     12,     0, ":::::*::::::::::"),
	(0,     0,     0,     ':',     2,     0, ":::::*::::::B:::"),
	(0,     0,     1,     ':',     2,     0, ":::::*::::::B:::"),
	(0,     0,     1,     'W',     4,     0, ":::::*::::::B:::"),
	(0,     0,     1,     '*',     5,     0, "::::W*::::::B:::"),
	(0,     0,     1,     'W',     13,     0, "::::W:::::::B:::"),
	(0,     0,     1,     ':',     13,     0, "::::W:::::::BW::"),
	(0,     0,     0,     '*',     9,     0, "::::W:::::::BW::"),
	(0,     0,     0,     'W',     12,     0, "::::W:::::::BW::"),
	(0,     0,     0,     '*',     6,     0, "::::W:::::::BW::"),
	(0,     0,     0,     'B',     9,     0, "::::W:::::::BW::"),
	(1,     1,     0,     'W',     13,     0, "::::W:::::::BW::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, "::::::::::::::B:"),
	(0,     0,     0,     'W',     7,     0, ":::::::::W::::B:"),
	(0,     0,     0,     'W',     13,     0, ":::::::::W::::B:"),
	(0,     0,     1,     '*',     13,     0, ":::::::::W::::B:"),
	(0,     0,     1,     '*',     10,     0, ":::::::::W:::*B:"),
	(0,     0,     0,     ':',     2,     0, ":::::::::W*::*B:"),
	(0,     0,     0,     '*',     13,     0, ":::::::::W*::*B:"),
	(0,     0,     1,     ':',     10,     0, ":::::::::W*::*B:"),
	(1,     0,     1,     'B',     8,     0, ":::::::::W*::*B:"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     4,     0, "::::::::::W::W::"),
	(0,     0,     0,     'B',     9,     0, "::::::::::W::W::"),
	(0,     0,     0,     'W',     5,     0, "::::::::::W::W::"),
	(0,     0,     0,     'B',     13,     0, "::::::::::W::W::"),
	(0,     0,     0,     'B',     7,     0, "::::::::::W::W::"),
	(0,     0,     1,     '*',     9,     0, "::::::::::W::W::"),
	(0,     0,     0,     'B',     6,     0, ":::::::::*W::W::"),
	(0,     0,     1,     'W',     13,     0, ":::::::::*W::W::"),
	(0,     0,     0,     ':',     7,     0, ":::::::::*W::W::"),
	(0,     0,     1,     '*',     9,     0, ":::::::::*W::W::"),
	(0,     1,     0,     ':',     6,     0, "::::::::::W::W::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     15,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":B::::::::::::::"),
	(0,     0,     1,     ':',     6,     0, ":B::::::::::::::"),
	(0,     1,     0,     '*',     2,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     1,     0, ":::::::::::::*::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::::::*::"),
	(0,     1,     0,     '*',     0,     0, "::::::::*::::*::"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     0, "::::::::::::::W:"),
	(0,     1,     0,     'B',     2,     0, "::::::::::::::W:"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, ":W::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "*W::::::::::::::"),
	(0,     0,     1,     '*',     2,     0, "*W::::::::::::::"),
	(0,     0,     1,     'W',     5,     0, "*W*:::::::::::::"),
	(0,     0,     1,     'W',     3,     0, "*W*::W::::::::::"),
	(0,     0,     0,     '*',     3,     0, "*W*W:W::::::::::"),
	(0,     0,     0,     'W',     10,     0, "*W*W:W::::::::::"),
	(0,     0,     0,     ':',     6,     0, "*W*W:W::::::::::"),
	(0,     0,     1,     ':',     14,     0, "*W*W:W::::::::::"),
	(0,     0,     1,     ':',     11,     0, "*W*W:W::::::::::"),
	(0,     0,     1,     'B',     0,     0, "*W*W:W::::::::::"),
	(0,     1,     0,     'B',     11,     0, "BW*W:W::::::::::"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     0,     0, ":::W:::::::::W::"),
	(0,     1,     0,     'B',     12,     0, ":::W:::::::::W::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, "::B:::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "::B:::::B:::::::"),
	(0,     0,     0,     ':',     10,     0, "::B:::::B:::::::"),
	(0,     0,     0,     'W',     3,     0, "::B:::::B:::::::"),
	(0,     0,     1,     ':',     8,     0, "::B:::::B:::::::"),
	(0,     0,     0,     '*',     0,     0, "::B:::::B:::::::"),
	(0,     1,     1,     'W',     12,     0, "::B:::::B:::::::"),
	(0,     0,     1,     '*',     1,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     3,     0, ":*::::::::::W:::"),
	(0,     1,     1,     '*',     5,     0, ":*:W::::::::W:::"),
	(0,     0,     1,     'W',     4,     0, ":::::*::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::::W*::::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::W*::::::::W:"),
	(0,     0,     0,     ':',     0,     0, "::*:W*::::::::W:"),
	(0,     0,     1,     'W',     5,     0, "::*:W*::::::::W:"),
	(0,     0,     1,     'B',     2,     0, "::*:WW::::::::W:"),
	(0,     0,     1,     ':',     0,     0, "::B:WW::::::::W:"),
	(0,     1,     0,     '*',     13,     0, "::B:WW::::::::W:"),
	(0,     1,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     11,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     11,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     9,     0, ":::::W::::::::::"),
	(0,     0,     1,     'B',     15,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     8,     0, ":::::W:::::::::B"),
	(0,     0,     0,     ':',     4,     0, ":::::W::W::::::B"),
	(0,     0,     1,     'W',     0,     0, ":::::W::W::::::B"),
	(0,     0,     1,     'W',     12,     0, "W::::W::W::::::B"),
	(0,     0,     0,     '*',     13,     0, "W::::W::W:::W::B"),
	(0,     0,     0,     'B',     1,     0, "W::::W::W:::W::B"),
	(0,     0,     0,     'B',     14,     0, "W::::W::W:::W::B"),
	(0,     1,     0,     '*',     13,     0, "W::::W::W:::W::B"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     15,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     6,     0, ":::::::::::B::::"),
	(0,     0,     0,     '*',     3,     0, ":::::::::::B::::"),
	(0,     0,     1,     'W',     10,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     13,     0, "::::::::::WB::::"),
	(0,     0,     1,     '*',     14,     0, "::::::::::WB::::"),
	(0,     0,     1,     'W',     8,     0, "::::::::::WB::*:"),
	(0,     0,     0,     'W',     7,     0, "::::::::W:WB::*:"),
	(0,     0,     1,     '*',     15,     0, "::::::::W:WB::*:"),
	(0,     0,     0,     'B',     1,     0, "::::::::W:WB::**"),
	(0,     0,     0,     '*',     12,     0, "::::::::W:WB::**"),
	(0,     0,     1,     ':',     2,     0, "::::::::W:WB::**"),
	(0,     0,     1,     'W',     12,     0, "::::::::W:WB::**"),
	(0,     0,     1,     '*',     6,     0, "::::::::W:WBW:**"),
	(1,     0,     0,     'W',     12,     0, "::::::*:W:WBW:**"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(1,     0,     1,     'W',     5,     0, ":W::::::::::::::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     3,     0, "::::::::::::W:::"),
	(0,     1,     0,     ':',     10,     0, ":::*::::::::W:::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::::::::::::B::"),
	(0,     0,     1,     'W',     7,     0, ":::::::::::::B::"),
	(0,     0,     1,     ':',     13,     0, ":::::::W:::::B::"),
	(0,     0,     1,     '*',     2,     0, ":::::::W:::::B::"),
	(0,     0,     1,     ':',     4,     0, "::*::::W:::::B::"),
	(0,     0,     0,     'B',     4,     0, "::*::::W:::::B::"),
	(0,     0,     0,     '*',     7,     0, "::*::::W:::::B::"),
	(0,     0,     0,     '*',     11,     0, "::*::::W:::::B::"),
	(0,     0,     0,     'W',     15,     0, "::*::::W:::::B::"),
	(0,     1,     1,     'B',     9,     0, "::*::::W:::::B::"),
	(0,     0,     1,     'B',     12,     0, ":::::::::B::::::"),
	(0,     0,     1,     'W',     4,     0, ":::::::::B::B:::"),
	(0,     0,     1,     'B',     9,     0, "::::W::::B::B:::"),
	(0,     0,     0,     ':',     1,     0, "::::W::::B::B:::"),
	(0,     0,     0,     'B',     12,     0, "::::W::::B::B:::"),
	(0,     0,     1,     'W',     2,     0, "::::W::::B::B:::"),
	(0,     0,     0,     'W',     7,     0, "::W:W::::B::B:::"),
	(0,     1,     1,     ':',     12,     0, "::W:W::::B::B:::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     0, ":W::::::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":W::::::::::::::"),
	(0,     0,     0,     'W',     10,     0, ":W::::W:::::::::"),
	(0,     0,     1,     ':',     3,     0, ":W::::W:::::::::"),
	(0,     0,     1,     'B',     2,     0, ":W::::W:::::::::"),
	(0,     0,     0,     '*',     13,     0, ":WB:::W:::::::::"),
	(0,     0,     0,     'B',     0,     0, ":WB:::W:::::::::"),
	(0,     0,     0,     '*',     10,     0, ":WB:::W:::::::::"),
	(0,     0,     1,     'W',     8,     0, ":WB:::W:::::::::"),
	(0,     0,     1,     '*',     8,     0, ":WB:::W:W:::::::"),
	(0,     0,     0,     'B',     4,     0, ":WB:::W:B:::::::"),
	(0,     0,     1,     ':',     12,     0, ":WB:::W:B:::::::"),
	(0,     0,     0,     'B',     8,     0, ":WB:::W:B:::::::"),
	(1,     0,     0,     'B',     4,     0, ":WB:::W:B:::::::"),
	(0,     1,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     8,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     12,     0, ":::*::::W:::::::"),
	(0,     0,     1,     'B',     3,     0, ":::*::::W:::::::"),
	(0,     1,     1,     'B',     10,     0, ":::B::::W:::::::"),
	(0,     1,     0,     'W',     12,     0, "::::::::::B:::::"),
	(0,     0,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::::::::::::*:"),
	(1,     1,     0,     '*',     4,     0, "::::::::::::::*:"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::B:::B::::::::"),
	(0,     0,     1,     'B',     0,     0, ":::B:::B::::::::"),
	(0,     0,     0,     ':',     3,     0, "B::B:::B::::::::"),
	(0,     0,     1,     ':',     6,     0, "B::B:::B::::::::"),
	(0,     0,     0,     'B',     5,     0, "B::B:::B::::::::"),
	(0,     0,     1,     ':',     1,     0, "B::B:::B::::::::"),
	(0,     0,     0,     'W',     12,     0, "B::B:::B::::::::"),
	(0,     0,     0,     'W',     3,     0, "B::B:::B::::::::"),
	(0,     0,     0,     '*',     7,     0, "B::B:::B::::::::"),
	(0,     0,     1,     'B',     0,     0, "B::B:::B::::::::"),
	(0,     0,     1,     'B',     15,     0, "B::B:::B::::::::"),
	(0,     0,     0,     ':',     5,     0, "B::B:::B:::::::B"),
	(0,     0,     1,     '*',     14,     0, "B::B:::B:::::::B"),
	(0,     0,     1,     '*',     11,     0, "B::B:::B::::::*B"),
	(0,     0,     1,     ':',     1,     0, "B::B:::B:::*::*B"),
	(0,     0,     1,     ':',     10,     0, "B::B:::B:::*::*B"),
	(0,     0,     1,     'B',     6,     0, "B::B:::B:::*::*B"),
	(0,     0,     0,     '*',     0,     0, "B::B::BB:::*::*B"),
	(0,     0,     0,     '*',     7,     0, "B::B::BB:::*::*B"),
	(0,     0,     0,     ':',     1,     0, "B::B::BB:::*::*B"),
	(0,     0,     1,     '*',     6,     0, "B::B::BB:::*::*B"),
	(0,     0,     0,     ':',     3,     0, "B::B::WB:::*::*B"),
	(0,     0,     1,     ':',     15,     0, "B::B::WB:::*::*B"),
	(0,     0,     1,     'B',     13,     0, "B::B::WB:::*::*B"),
	(0,     0,     1,     'W',     9,     0, "B::B::WB:::*:B*B"),
	(0,     0,     0,     'W',     6,     0, "B::B::WB:W:*:B*B"),
	(0,     0,     0,     'B',     3,     0, "B::B::WB:W:*:B*B"),
	(0,     1,     0,     ':',     4,     0, "B::B::WB:W:*:B*B"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":W::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, ":B::::::::::::::"),
	(0,     1,     1,     ':',     13,     0, ":B::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     15,     0, ":::::::::::::B::"),
	(0,     0,     1,     ':',     11,     0, ":::::::::::::::B"),
	(0,     0,     0,     'B',     6,     0, ":::::::::::::::B"),
	(0,     0,     1,     'B',     6,     0, ":::::::::::::::B"),
	(0,     0,     0,     'B',     0,     0, "::::::B::::::::B"),
	(0,     1,     1,     ':',     13,     0, "::::::B::::::::B"),
	(0,     0,     0,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     0, "*:::::::::::::::"),
	(0,     0,     1,     ':',     0,     0, "*::::::::B::::::"),
	(0,     0,     0,     'B',     10,     0, "*::::::::B::::::"),
	(0,     0,     0,     'W',     3,     0, "*::::::::B::::::"),
	(0,     0,     1,     'W',     7,     0, "*::::::::B::::::"),
	(0,     0,     0,     'W',     1,     0, "*::::::W:B::::::"),
	(0,     0,     0,     'W',     15,     0, "*::::::W:B::::::"),
	(0,     0,     0,     ':',     8,     0, "*::::::W:B::::::"),
	(0,     0,     1,     'W',     7,     0, "*::::::W:B::::::"),
	(0,     0,     1,     '*',     13,     0, "*::::::W:B::::::"),
	(0,     0,     0,     'B',     1,     0, "*::::::W:B:::*::"),
	(0,     0,     1,     'W',     6,     0, "*::::::W:B:::*::"),
	(0,     0,     0,     'B',     15,     0, "*:::::WW:B:::*::"),
	(0,     0,     1,     'W',     10,     0, "*:::::WW:B:::*::"),
	(0,     0,     1,     'B',     4,     0, "*:::::WW:BW::*::"),
	(0,     0,     0,     'B',     13,     0, "*:::B:WW:BW::*::"),
	(0,     0,     1,     ':',     5,     0, "*:::B:WW:BW::*::"),
	(0,     0,     0,     'B',     1,     0, "*:::B:WW:BW::*::"),
	(0,     0,     1,     'B',     8,     0, "*:::B:WW:BW::*::"),
	(0,     0,     0,     'W',     14,     0, "*:::B:WWBBW::*::"),
	(0,     0,     0,     'B',     9,     0, "*:::B:WWBBW::*::"),
	(0,     0,     0,     'W',     0,     0, "*:::B:WWBBW::*::"),
	(0,     0,     1,     'B',     11,     0, "*:::B:WWBBW::*::"),
	(0,     0,     0,     ':',     8,     0, "*:::B:WWBBWB:*::"),
	(0,     0,     0,     ':',     9,     0, "*:::B:WWBBWB:*::"),
	(0,     0,     1,     '*',     15,     0, "*:::B:WWBBWB:*::"),
	(0,     0,     1,     'B',     10,     0, "*:::B:WWBBWB:*:*"),
	(0,     0,     1,     'W',     3,     0, "*:::B:WWBBBB:*:*"),
	(0,     0,     0,     'W',     6,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     1,     ':',     6,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     0,     'W',     5,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     1,     'B',     9,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     0,     'W',     5,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     0,     ':',     15,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     1,     'B',     5,     0, "*::WB:WWBBBB:*:*"),
	(0,     0,     0,     ':',     15,     0, "*::WBBWWBBBB:*:*"),
	(0,     0,     1,     ':',     10,     0, "*::WBBWWBBBB:*:*"),
	(0,     0,     1,     'B',     3,     0, "*::WBBWWBBBB:*:*"),
	(0,     0,     0,     ':',     10,     0, "*::BBBWWBBBB:*:*"),
	(0,     0,     1,     ':',     5,     0, "*::BBBWWBBBB:*:*"),
	(0,     0,     1,     '*',     1,     0, "*::BBBWWBBBB:*:*"),
	(0,     0,     0,     ':',     3,     0, "**:BBBWWBBBB:*:*"),
	(0,     0,     0,     'W',     4,     0, "**:BBBWWBBBB:*:*"),
	(0,     0,     0,     '*',     2,     0, "**:BBBWWBBBB:*:*"),
	(0,     0,     1,     'W',     8,     0, "**:BBBWWBBBB:*:*"),
	(0,     0,     0,     ':',     10,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     0,     'W',     3,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     0,     ':',     4,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     0,     'B',     3,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     0,     ':',     9,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     0,     'B',     9,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     1,     ':',     14,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     1,     'W',     2,     0, "**:BBBWWWBBB:*:*"),
	(0,     0,     0,     'B',     8,     0, "**WBBBWWWBBB:*:*"),
	(0,     0,     1,     'W',     15,     0, "**WBBBWWWBBB:*:*"),
	(0,     1,     1,     'W',     0,     0, "**WBBBWWWBBB:*:W"),
	(0,     0,     0,     ':',     12,     0, "W:::::::::::::::"),
	(0,     0,     0,     ':',     1,     0, "W:::::::::::::::"),
	(0,     0,     0,     'W',     7,     0, "W:::::::::::::::"),
	(0,     1,     1,     ':',     11,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, ":*::::::::B:::::"),
	(0,     0,     0,     '*',     12,     0, ":*::W:::::B:::::"),
	(0,     0,     0,     ':',     4,     0, ":*::W:::::B:::::"),
	(0,     0,     1,     'B',     11,     0, ":*::W:::::B:::::"),
	(0,     0,     1,     'B',     11,     0, ":*::W:::::BB::::"),
	(0,     0,     1,     '*',     12,     0, ":*::W:::::BB::::"),
	(0,     0,     1,     'B',     8,     0, ":*::W:::::BB*:::"),
	(0,     0,     1,     '*',     9,     0, ":*::W:::B:BB*:::"),
	(0,     1,     1,     'W',     5,     0, ":*::W:::B*BB*:::"),
	(0,     0,     0,     ':',     10,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     9,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     7,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     12,     0, ":::::W:W::::::::"),
	(0,     1,     0,     '*',     5,     0, ":::::W:W::::::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     13,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::::::::::::B:"),
	(0,     1,     1,     'W',     9,     0, "::::::::::::::B:"),
	(0,     0,     1,     '*',     11,     0, ":::::::::W::::::"),
	(0,     0,     0,     'W',     2,     0, ":::::::::W:*::::"),
	(0,     0,     1,     'W',     2,     0, ":::::::::W:*::::"),
	(0,     0,     1,     ':',     6,     0, "::W::::::W:*::::"),
	(0,     0,     0,     'B',     4,     0, "::W::::::W:*::::"),
	(0,     0,     1,     'W',     4,     0, "::W::::::W:*::::"),
	(0,     0,     1,     '*',     13,     0, "::W:W::::W:*::::"),
	(0,     0,     1,     'W',     1,     0, "::W:W::::W:*:*::"),
	(0,     0,     1,     ':',     14,     0, ":WW:W::::W:*:*::"),
	(0,     0,     0,     'B',     1,     0, ":WW:W::::W:*:*::"),
	(0,     0,     1,     '*',     12,     0, ":WW:W::::W:*:*::"),
	(0,     0,     0,     ':',     4,     0, ":WW:W::::W:***::"),
	(0,     0,     0,     'W',     12,     0, ":WW:W::::W:***::"),
	(0,     1,     0,     '*',     3,     0, ":WW:W::::W:***::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     10,     0, ":B::::::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":B::::::::::::::"),
	(0,     0,     0,     ':',     14,     0, ":B::::::::::::::"),
	(0,     0,     1,     'B',     5,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":B:::B::::::::::"),
	(0,     0,     0,     'B',     0,     0, ":W:::B::::::::::"),
	(0,     1,     0,     '*',     15,     0, ":W:::B::::::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, "::::B:::::::::::"),
	(0,     0,     0,     'W',     12,     0, "::::B:::::::::::"),
	(0,     0,     0,     ':',     9,     0, "::::B:::::::::::"),
	(0,     0,     0,     ':',     0,     0, "::::B:::::::::::"),
	(0,     0,     0,     '*',     1,     0, "::::B:::::::::::"),
	(0,     1,     1,     '*',     4,     0, "::::B:::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::::*:::::::::::"),
	(0,     0,     0,     ':',     9,     0, "::::*:::::::::::"),
	(0,     0,     1,     'B',     2,     0, "::::*:::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::B:*:::::::::::"),
	(0,     0,     0,     '*',     5,     0, "::B:*:::::::::::"),
	(0,     0,     1,     'B',     5,     0, "::B:*:::::::::::"),
	(0,     0,     1,     'W',     8,     0, "::B:*B::::::::::"),
	(0,     0,     0,     'B',     7,     0, "::B:*B::W:::::::"),
	(0,     0,     1,     'W',     11,     0, "::B:*B::W:::::::"),
	(0,     0,     1,     'B',     7,     0, "::B:*B::W::W::::"),
	(0,     0,     1,     'B',     0,     0, "::B:*B:BW::W::::"),
	(0,     0,     1,     ':',     12,     0, "B:B:*B:BW::W::::"),
	(0,     1,     1,     'W',     10,     0, "B:B:*B:BW::W::::"),
	(0,     0,     1,     '*',     14,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     3,     0, "::::::::::W:::*:"),
	(0,     0,     0,     'W',     5,     0, "::::::::::W:::*:"),
	(0,     0,     0,     '*',     12,     0, "::::::::::W:::*:"),
	(0,     0,     1,     'B',     2,     0, "::::::::::W:::*:"),
	(0,     0,     1,     'W',     9,     0, "::B:::::::W:::*:"),
	(0,     0,     1,     ':',     10,     0, "::B::::::WW:::*:"),
	(0,     0,     0,     'B',     15,     0, "::B::::::WW:::*:"),
	(0,     0,     1,     'W',     6,     0, "::B::::::WW:::*:"),
	(0,     0,     1,     ':',     14,     0, "::B:::W::WW:::*:"),
	(0,     0,     1,     'W',     4,     0, "::B:::W::WW:::*:"),
	(0,     0,     0,     'B',     14,     0, "::B:W:W::WW:::*:"),
	(0,     0,     1,     'W',     14,     0, "::B:W:W::WW:::*:"),
	(0,     0,     1,     'W',     3,     0, "::B:W:W::WW:::W:"),
	(0,     0,     1,     '*',     0,     0, "::BWW:W::WW:::W:"),
	(0,     0,     0,     ':',     11,     0, "*:BWW:W::WW:::W:"),
	(0,     0,     1,     ':',     15,     0, "*:BWW:W::WW:::W:"),
	(0,     0,     1,     'W',     14,     0, "*:BWW:W::WW:::W:"),
	(0,     0,     0,     ':',     3,     0, "*:BWW:W::WW:::W:"),
	(0,     0,     1,     'W',     1,     0, "*:BWW:W::WW:::W:"),
	(0,     0,     0,     '*',     13,     0, "*WBWW:W::WW:::W:"),
	(0,     0,     1,     'W',     4,     0, "*WBWW:W::WW:::W:"),
	(0,     0,     0,     'B',     13,     0, "*WBWW:W::WW:::W:"),
	(0,     0,     1,     'B',     11,     0, "*WBWW:W::WW:::W:"),
	(0,     0,     0,     '*',     13,     0, "*WBWW:W::WWB::W:"),
	(0,     0,     1,     'W',     15,     0, "*WBWW:W::WWB::W:"),
	(0,     0,     0,     ':',     13,     0, "*WBWW:W::WWB::WW"),
	(0,     0,     0,     'W',     8,     0, "*WBWW:W::WWB::WW"),
	(0,     0,     0,     'B',     10,     0, "*WBWW:W::WWB::WW"),
	(0,     0,     1,     'W',     8,     0, "*WBWW:W::WWB::WW"),
	(0,     0,     1,     'B',     8,     0, "*WBWW:W:WWWB::WW"),
	(0,     0,     0,     ':',     15,     0, "*WBWW:W:BWWB::WW"),
	(0,     0,     0,     '*',     1,     0, "*WBWW:W:BWWB::WW"),
	(0,     0,     0,     ':',     14,     0, "*WBWW:W:BWWB::WW"),
	(0,     0,     1,     ':',     12,     0, "*WBWW:W:BWWB::WW"),
	(0,     1,     1,     '*',     4,     0, "*WBWW:W:BWWB::WW"),
	(0,     0,     1,     'W',     5,     0, "::::*:::::::::::"),
	(0,     0,     0,     '*',     8,     0, "::::*W::::::::::"),
	(0,     0,     1,     'W',     15,     0, "::::*W::::::::::"),
	(0,     0,     1,     '*',     11,     0, "::::*W:::::::::W"),
	(0,     0,     1,     'B',     5,     0, "::::*W:::::*:::W"),
	(0,     1,     0,     'B',     11,     0, "::::*B:::::*:::W"),
	(0,     1,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::::::::B:::::"),
	(0,     0,     0,     'B',     1,     0, "::::::::::B:::::"),
	(0,     0,     0,     'B',     8,     0, "::::::::::B:::::"),
	(0,     1,     1,     'W',     6,     0, "::::::::::B:::::"),
	(0,     0,     0,     'W',     0,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     10,     0, "::::::W:::::::::"),
	(0,     0,     1,     ':',     3,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     3,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     12,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     11,     0, "::::::W:::::B:::"),
	(0,     0,     0,     '*',     2,     0, "::::::W:::::B:::"),
	(0,     0,     1,     ':',     4,     0, "::::::W:::::B:::"),
	(0,     0,     0,     'W',     14,     0, "::::::W:::::B:::"),
	(0,     0,     1,     'B',     13,     0, "::::::W:::::B:::"),
	(0,     0,     1,     '*',     9,     0, "::::::W:::::BB::"),
	(0,     0,     0,     '*',     13,     0, "::::::W::*::BB::"),
	(0,     0,     0,     ':',     11,     0, "::::::W::*::BB::"),
	(0,     0,     0,     ':',     11,     0, "::::::W::*::BB::"),
	(0,     0,     1,     'W',     14,     0, "::::::W::*::BB::"),
	(0,     0,     0,     'B',     13,     0, "::::::W::*::BBW:"),
	(0,     1,     1,     'B',     8,     0, "::::::W::*::BBW:"),
	(0,     0,     0,     'B',     8,     0, "::::::::B:::::::"),
	(0,     0,     0,     '*',     14,     0, "::::::::B:::::::"),
	(0,     0,     1,     'B',     13,     0, "::::::::B:::::::"),
	(0,     0,     0,     'B',     1,     0, "::::::::B::::B::"),
	(0,     0,     1,     'W',     4,     0, "::::::::B::::B::"),
	(0,     0,     1,     'B',     15,     0, "::::W:::B::::B::"),
	(0,     0,     1,     'B',     15,     0, "::::W:::B::::B:B"),
	(0,     1,     0,     'W',     12,     0, "::::W:::B::::B:B"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     8,     0, ":::::::::::::::*"),
	(0,     0,     0,     'W',     5,     0, ":::::::::::::::*"),
	(0,     0,     1,     ':',     0,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     1,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     4,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     14,     0, ":::::::::::::::*"),
	(0,     0,     1,     ':',     7,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     1,     0, ":::::::::::::::*"),
	(0,     0,     0,     ':',     9,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     10,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     0,     0, ":::::::::::::::*"),
	(0,     0,     0,     'B',     7,     0, ":::::::::::::::*"),
	(0,     1,     0,     '*',     12,     0, ":::::::::::::::*"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::::W::::::::::"),
	(0,     0,     0,     'B',     9,     0, ":::::W:::::::W::"),
	(0,     0,     0,     'W',     8,     0, ":::::W:::::::W::"),
	(0,     0,     0,     'B',     10,     0, ":::::W:::::::W::"),
	(0,     0,     1,     '*',     6,     0, ":::::W:::::::W::"),
	(0,     0,     1,     ':',     13,     0, ":::::W*::::::W::"),
	(0,     0,     1,     'B',     8,     0, ":::::W*::::::W::"),
	(0,     0,     0,     ':',     8,     0, ":::::W*:B::::W::"),
	(0,     0,     1,     'B',     6,     0, ":::::W*:B::::W::"),
	(0,     0,     0,     ':',     10,     0, ":::::WB:B::::W::"),
	(0,     0,     0,     'W',     5,     0, ":::::WB:B::::W::"),
	(0,     0,     0,     'B',     12,     0, ":::::WB:B::::W::"),
	(0,     1,     1,     'B',     5,     0, ":::::WB:B::::W::"),
	(0,     0,     1,     '*',     11,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     14,     0, ":::::B:::::*::::"),
	(0,     0,     1,     'B',     12,     0, ":::::B:::::*::*:"),
	(0,     1,     1,     'W',     3,     0, ":::::B:::::*B:*:"),
	(0,     0,     0,     ':',     14,     0, ":::W::::::::::::"),
	(0,     0,     1,     '*',     5,     0, ":::W::::::::::::"),
	(0,     0,     0,     'W',     8,     0, ":::W:*::::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::W:*::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":::W:*::::::::::"),
	(0,     0,     0,     ':',     1,     0, ":::W:*W:::::::::"),
	(0,     0,     0,     'W',     0,     0, ":::W:*W:::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::W:*W:::::::::"),
	(0,     0,     1,     'B',     10,     0, ":::W:*W:::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::W:*W:::B:::::"),
	(0,     0,     0,     'B',     10,     0, ":::W:*W:::B:::::"),
	(0,     0,     0,     'B',     7,     0, ":::W:*W:::B:::::"),
	(0,     0,     0,     ':',     12,     0, ":::W:*W:::B:::::"),
	(0,     0,     1,     '*',     5,     0, ":::W:*W:::B:::::"),
	(0,     0,     1,     ':',     13,     0, ":::W::W:::B:::::"),
	(0,     0,     1,     'W',     6,     0, ":::W::W:::B:::::"),
	(0,     0,     1,     '*',     12,     0, ":::W::W:::B:::::"),
	(0,     0,     0,     ':',     13,     0, ":::W::W:::B:*:::"),
	(0,     0,     0,     'B',     4,     0, ":::W::W:::B:*:::"),
	(0,     0,     0,     'W',     0,     0, ":::W::W:::B:*:::"),
	(0,     0,     1,     'B',     5,     0, ":::W::W:::B:*:::"),
	(0,     0,     0,     ':',     6,     0, ":::W:BW:::B:*:::"),
	(0,     0,     0,     'B',     6,     0, ":::W:BW:::B:*:::"),
	(0,     0,     1,     'W',     9,     0, ":::W:BW:::B:*:::"),
	(0,     0,     0,     'B',     14,     0, ":::W:BW::WB:*:::"),
	(0,     0,     0,     ':',     4,     0, ":::W:BW::WB:*:::"),
	(0,     0,     1,     'W',     8,     0, ":::W:BW::WB:*:::"),
	(0,     0,     1,     'B',     11,     0, ":::W:BW:WWB:*:::"),
	(0,     0,     0,     '*',     11,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     0,     ':',     9,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     0,     'B',     10,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     1,     'B',     5,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     0,     'B',     14,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     0,     '*',     6,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     1,     'B',     11,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     0,     'W',     1,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     1,     'W',     15,     0, ":::W:BW:WWBB*:::"),
	(0,     0,     1,     'W',     1,     0, ":::W:BW:WWBB*::W"),
	(0,     0,     0,     'B',     15,     0, ":W:W:BW:WWBB*::W"),
	(0,     0,     1,     'B',     3,     0, ":W:W:BW:WWBB*::W"),
	(0,     0,     1,     ':',     15,     0, ":W:B:BW:WWBB*::W"),
	(0,     0,     1,     ':',     6,     0, ":W:B:BW:WWBB*::W"),
	(0,     0,     0,     'B',     0,     0, ":W:B:BW:WWBB*::W"),
	(0,     0,     0,     ':',     1,     0, ":W:B:BW:WWBB*::W"),
	(0,     0,     1,     'B',     8,     0, ":W:B:BW:WWBB*::W"),
	(0,     0,     0,     ':',     1,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     0,     ':',     13,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     0,     'W',     10,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     1,     ':',     13,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     0,     '*',     4,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     0,     '*',     10,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     1,     ':',     8,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     0,     'B',     0,     0, ":W:B:BW:BWBB*::W"),
	(0,     0,     0,     'W',     9,     0, ":W:B:BW:BWBB*::W"),
	(0,     1,     1,     ':',     2,     0, ":W:B:BW:BWBB*::W"),
	(0,     1,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "::::::::::::B:::"),
	(0,     0,     1,     '*',     14,     0, "::::::::::::B:::"),
	(0,     0,     0,     ':',     6,     0, "::::::::::::B:*:"),
	(0,     0,     1,     ':',     13,     0, "::::::::::::B:*:"),
	(0,     0,     0,     '*',     14,     0, "::::::::::::B:*:"),
	(0,     0,     1,     'B',     4,     0, "::::::::::::B:*:"),
	(0,     0,     1,     ':',     7,     0, "::::B:::::::B:*:"),
	(0,     0,     1,     'W',     12,     0, "::::B:::::::B:*:"),
	(0,     0,     0,     'B',     11,     0, "::::B:::::::W:*:"),
	(0,     0,     1,     ':',     8,     0, "::::B:::::::W:*:"),
	(0,     0,     0,     'B',     9,     0, "::::B:::::::W:*:"),
	(0,     0,     1,     '*',     0,     0, "::::B:::::::W:*:"),
	(0,     0,     0,     'W',     14,     0, "*:::B:::::::W:*:"),
	(0,     0,     0,     '*',     6,     0, "*:::B:::::::W:*:"),
	(0,     0,     1,     'B',     1,     0, "*:::B:::::::W:*:"),
	(0,     0,     0,     '*',     11,     0, "*B::B:::::::W:*:"),
	(0,     0,     0,     'W',     4,     0, "*B::B:::::::W:*:"),
	(0,     0,     0,     'B',     4,     0, "*B::B:::::::W:*:"),
	(0,     0,     0,     'B',     10,     0, "*B::B:::::::W:*:"),
	(0,     0,     1,     '*',     1,     0, "*B::B:::::::W:*:"),
	(0,     0,     1,     '*',     6,     0, "*W::B:::::::W:*:"),
	(0,     0,     1,     ':',     8,     0, "*W::B:*:::::W:*:"),
	(0,     0,     1,     ':',     0,     0, "*W::B:*:::::W:*:"),
	(0,     0,     0,     'B',     11,     0, "*W::B:*:::::W:*:"),
	(0,     0,     1,     'B',     13,     0, "*W::B:*:::::W:*:"),
	(0,     0,     0,     '*',     11,     0, "*W::B:*:::::WB*:"),
	(0,     0,     1,     'W',     9,     0, "*W::B:*:::::WB*:"),
	(0,     0,     0,     ':',     15,     0, "*W::B:*::W::WB*:"),
	(0,     0,     1,     'W',     1,     0, "*W::B:*::W::WB*:"),
	(0,     0,     0,     'W',     8,     0, "*W::B:*::W::WB*:"),
	(0,     0,     0,     'B',     7,     0, "*W::B:*::W::WB*:"),
	(0,     0,     1,     '*',     12,     0, "*W::B:*::W::WB*:"),
	(0,     0,     1,     '*',     9,     0, "*W::B:*::W::BB*:"),
	(0,     0,     1,     'W',     3,     0, "*W::B:*::B::BB*:"),
	(0,     0,     0,     ':',     12,     0, "*W:WB:*::B::BB*:"),
	(0,     0,     0,     '*',     9,     0, "*W:WB:*::B::BB*:"),
	(0,     0,     1,     '*',     9,     0, "*W:WB:*::B::BB*:"),
	(0,     0,     1,     '*',     5,     0, "*W:WB:*::W::BB*:"),
	(0,     0,     0,     'B',     5,     0, "*W:WB**::W::BB*:"),
	(0,     0,     1,     '*',     11,     0, "*W:WB**::W::BB*:"),
	(0,     0,     0,     'B',     13,     0, "*W:WB**::W:*BB*:"),
	(0,     0,     0,     '*',     3,     0, "*W:WB**::W:*BB*:"),
	(0,     0,     1,     'B',     10,     0, "*W:WB**::W:*BB*:"),
	(0,     0,     0,     'W',     11,     0, "*W:WB**::WB*BB*:"),
	(0,     0,     0,     'B',     9,     0, "*W:WB**::WB*BB*:"),
	(0,     0,     0,     'W',     9,     0, "*W:WB**::WB*BB*:"),
	(0,     0,     0,     ':',     7,     0, "*W:WB**::WB*BB*:"),
	(0,     0,     0,     ':',     10,     0, "*W:WB**::WB*BB*:"),
	(0,     1,     1,     'W',     8,     0, "*W:WB**::WB*BB*:"),
	(0,     0,     0,     'B',     15,     0, "::::::::W:::::::"),
	(0,     0,     0,     'W',     15,     0, "::::::::W:::::::"),
	(0,     0,     0,     'B',     7,     0, "::::::::W:::::::"),
	(0,     0,     1,     'B',     2,     0, "::::::::W:::::::"),
	(0,     1,     1,     '*',     4,     0, "::B:::::W:::::::"),
	(0,     0,     1,     '*',     5,     0, "::::*:::::::::::"),
	(0,     0,     1,     'B',     11,     0, "::::**::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::::**:::::B::::"),
	(0,     0,     0,     ':',     15,     0, "::::**:::::B::::"),
	(0,     0,     0,     'B',     9,     0, "::::**:::::B::::"),
	(0,     0,     1,     'W',     3,     0, "::::**:::::B::::"),
	(0,     0,     1,     ':',     6,     0, ":::W**:::::B::::"),
	(0,     0,     1,     'B',     7,     0, ":::W**:::::B::::"),
	(0,     0,     1,     '*',     12,     0, ":::W**:B:::B::::"),
	(0,     0,     0,     'B',     9,     0, ":::W**:B:::B*:::"),
	(0,     0,     0,     'W',     2,     0, ":::W**:B:::B*:::"),
	(0,     0,     1,     'B',     9,     0, ":::W**:B:::B*:::"),
	(0,     0,     1,     'B',     2,     0, ":::W**:B:B:B*:::"),
	(0,     0,     0,     '*',     12,     0, "::BW**:B:B:B*:::"),
	(0,     0,     0,     '*',     2,     0, "::BW**:B:B:B*:::"),
	(0,     0,     0,     'B',     14,     0, "::BW**:B:B:B*:::"),
	(0,     0,     1,     ':',     11,     0, "::BW**:B:B:B*:::"),
	(0,     0,     0,     '*',     14,     0, "::BW**:B:B:B*:::"),
	(0,     0,     1,     '*',     15,     0, "::BW**:B:B:B*:::"),
	(0,     0,     1,     'B',     1,     0, "::BW**:B:B:B*::*"),
	(0,     1,     1,     '*',     12,     0, ":BBW**:B:B:B*::*"),
	(0,     0,     0,     ':',     14,     0, "::::::::::::*:::"),
	(0,     0,     0,     'B',     5,     0, "::::::::::::*:::"),
	(0,     1,     0,     '*',     3,     0, "::::::::::::*:::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     11,     0, ":::::::::::B::::"),
	(0,     0,     1,     ':',     11,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     9,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     2,     0, ":::::::::*:B::::"),
	(0,     0,     0,     'W',     5,     0, "::*::::::*:B::::"),
	(0,     0,     0,     'B',     12,     0, "::*::::::*:B::::"),
	(0,     0,     1,     'W',     2,     0, "::*::::::*:B::::"),
	(1,     0,     0,     ':',     6,     0, "::W::::::*:B::::"),
	(0,     1,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     0, "::::::::W:::::::"),
	(0,     0,     0,     'W',     11,     0, "W:::::::W:::::::"),
	(0,     0,     0,     '*',     9,     0, "W:::::::W:::::::"),
	(0,     0,     0,     '*',     9,     0, "W:::::::W:::::::"),
	(0,     0,     1,     '*',     14,     0, "W:::::::W:::::::"),
	(0,     1,     1,     '*',     8,     0, "W:::::::W:::::*:"),
	(0,     0,     0,     ':',     7,     0, "::::::::*:::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::::*:::::::"),
	(0,     0,     0,     ':',     2,     0, "::::::::*:::::::"),
	(0,     0,     0,     '*',     7,     0, "::::::::*:::::::"),
	(0,     0,     0,     '*',     15,     0, "::::::::*:::::::"),
	(0,     0,     1,     ':',     0,     0, "::::::::*:::::::"),
	(0,     0,     0,     'B',     13,     0, "::::::::*:::::::"),
	(0,     0,     0,     'B',     1,     0, "::::::::*:::::::"),
	(0,     0,     0,     'W',     7,     0, "::::::::*:::::::"),
	(0,     1,     0,     'B',     6,     0, "::::::::*:::::::"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     0, "*:::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     14,     0, "*::::::::::B::::"),
	(0,     0,     0,     '*',     14,     0, "*::::::::::B::::"),
	(0,     1,     1,     ':',     3,     0, "*::::::::::B::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     8,     0, "B:::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, "B:::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "B:::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, "B:::::::::::::::"),
	(1,     0,     0,     ':',     3,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     3,     1, "::::::::::::::::"),
	(1,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, "::::B:::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::B:::::::::::"),
	(0,     0,     1,     '*',     6,     0, "::::B:::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::B:*:::::::::"),
	(0,     0,     1,     '*',     13,     0, "::::B:*:::::::::"),
	(0,     0,     1,     '*',     5,     0, "::::B:*::::::*::"),
	(0,     1,     0,     'W',     1,     0, "::::B**::::::*::"),
	(0,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, ":W::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, ":W::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, ":W::::::B:::::::"),
	(0,     1,     1,     'W',     12,     0, ":W::::::B:::::::"),
	(0,     0,     0,     ':',     1,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     3,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     1,     0, "::::::::::::W:::"),
	(0,     0,     1,     'B',     9,     0, ":W::::::::::W:::"),
	(0,     0,     0,     ':',     0,     0, ":W:::::::B::W:::"),
	(0,     0,     0,     'W',     7,     0, ":W:::::::B::W:::"),
	(0,     0,     0,     ':',     8,     0, ":W:::::::B::W:::"),
	(0,     1,     1,     'W',     2,     0, ":W:::::::B::W:::"),
	(0,     0,     1,     ':',     9,     0, "::W:::::::::::::"),
	(0,     0,     1,     ':',     10,     0, "::W:::::::::::::"),
	(0,     0,     0,     'W',     7,     0, "::W:::::::::::::"),
	(0,     0,     1,     'B',     4,     0, "::W:::::::::::::"),
	(0,     0,     1,     'B',     5,     0, "::W:B:::::::::::"),
	(0,     0,     1,     'B',     14,     0, "::W:BB::::::::::"),
	(0,     0,     0,     'W',     4,     0, "::W:BB::::::::B:"),
	(0,     0,     0,     ':',     5,     0, "::W:BB::::::::B:"),
	(0,     0,     1,     ':',     14,     0, "::W:BB::::::::B:"),
	(0,     0,     1,     'B',     11,     0, "::W:BB::::::::B:"),
	(0,     0,     1,     'B',     12,     0, "::W:BB:::::B::B:"),
	(0,     0,     0,     ':',     14,     0, "::W:BB:::::BB:B:"),
	(0,     0,     0,     '*',     15,     0, "::W:BB:::::BB:B:"),
	(0,     0,     0,     'B',     9,     0, "::W:BB:::::BB:B:"),
	(0,     0,     1,     '*',     1,     0, "::W:BB:::::BB:B:"),
	(0,     0,     1,     'W',     4,     0, ":*W:BB:::::BB:B:"),
	(0,     0,     1,     'W',     4,     0, ":*W:WB:::::BB:B:"),
	(0,     1,     0,     ':',     5,     0, ":*W:WB:::::BB:B:"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, ":::::::W::::::::"),
	(0,     0,     1,     '*',     0,     0, ":::B:::W::::::::"),
	(0,     1,     0,     '*',     2,     0, "*::B:::W::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::::::W::::::"),
	(0,     0,     1,     ':',     14,     0, ":::::::::W::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::::::W::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::W::::::"),
	(0,     0,     1,     'W',     12,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     15,     0, ":::::::::W::W:::"),
	(0,     1,     0,     '*',     10,     0, ":::::::::W::W:::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "::::::::B:::::::"),
	(0,     0,     1,     ':',     8,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     9,     0, "::::::::B:::::::"),
	(0,     0,     0,     '*',     7,     0, "::::::::B:::::::"),
	(0,     1,     1,     ':',     5,     0, "::::::::B:::::::"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, "B:::::::::::::::"),
	(0,     0,     1,     'W',     1,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     8,     0, "BW::::::::::::::"),
	(0,     0,     1,     '*',     10,     0, "BW::::::::::::::"),
	(0,     0,     1,     'B',     5,     0, "BW::::::::*:::::"),
	(0,     0,     1,     'B',     4,     0, "BW:::B::::*:::::"),
	(0,     1,     0,     'B',     6,     0, "BW::BB::::*:::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(1,     1,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     10,     0, "W:::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, "W:::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, "B:::::::::::::::"),
	(0,     0,     0,     'W',     6,     0, "B::B::::::::::::"),
	(0,     0,     0,     'B',     4,     0, "B::B::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "B::B::::::::::::"),
	(0,     0,     0,     ':',     7,     0, "B::B::::::::::::"),
	(0,     0,     1,     'B',     0,     0, "B::B::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "B::B::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "B::B::::::::::::"),
	(0,     0,     0,     'B',     3,     0, "B::BW:::::::::::"),
	(0,     0,     1,     '*',     7,     0, "B::BW:::::::::::"),
	(0,     0,     1,     ':',     9,     0, "B::BW::*::::::::"),
	(0,     0,     0,     'W',     9,     0, "B::BW::*::::::::"),
	(0,     0,     0,     'W',     0,     0, "B::BW::*::::::::"),
	(0,     0,     0,     ':',     7,     0, "B::BW::*::::::::"),
	(0,     0,     1,     ':',     12,     0, "B::BW::*::::::::"),
	(0,     0,     1,     'B',     3,     0, "B::BW::*::::::::"),
	(0,     0,     1,     ':',     8,     0, "B::BW::*::::::::"),
	(0,     0,     0,     'W',     11,     0, "B::BW::*::::::::"),
	(0,     0,     1,     ':',     3,     0, "B::BW::*::::::::"),
	(0,     0,     1,     'W',     5,     0, "B::BW::*::::::::"),
	(0,     0,     1,     'B',     6,     0, "B::BWW:*::::::::"),
	(0,     0,     1,     'W',     1,     0, "B::BWWB*::::::::"),
	(0,     0,     1,     'W',     13,     0, "BW:BWWB*::::::::"),
	(0,     0,     1,     '*',     8,     0, "BW:BWWB*:::::W::"),
	(0,     0,     1,     ':',     10,     0, "BW:BWWB**::::W::"),
	(0,     0,     1,     'B',     13,     0, "BW:BWWB**::::W::"),
	(0,     0,     0,     '*',     10,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     '*',     12,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     ':',     10,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     '*',     9,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     'W',     10,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     'W',     3,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     'W',     13,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     'B',     12,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     'W',     8,     0, "BW:BWWB**::::B::"),
	(0,     0,     1,     '*',     6,     0, "BW:BWWB**::::B::"),
	(0,     0,     0,     'W',     9,     0, "BW:BWWW**::::B::"),
	(0,     0,     1,     'W',     6,     0, "BW:BWWW**::::B::"),
	(0,     0,     0,     'B',     0,     0, "BW:BWWW**::::B::"),
	(0,     1,     0,     'W',     13,     0, "BW:BWWW**::::B::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::::::::::*::::"),
	(0,     0,     1,     '*',     1,     0, ":::::::::::*::::"),
	(0,     1,     1,     'B',     14,     0, ":*:::::::::*::::"),
	(0,     0,     0,     ':',     13,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     12,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     7,     0, "::::::::::::W:B:"),
	(0,     0,     0,     ':',     0,     0, ":::::::W::::W:B:"),
	(0,     0,     1,     'W',     3,     0, ":::::::W::::W:B:"),
	(0,     1,     0,     ':',     10,     0, ":::W:::W::::W:B:"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":*::::::::::::::"),
	(0,     0,     0,     ':',     1,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     6,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, ":*::::B:::::::::"),
	(0,     0,     1,     'W',     13,     0, ":*:B::B:::::::::"),
	(0,     0,     0,     ':',     4,     0, ":*:B::B::::::W::"),
	(0,     0,     0,     ':',     3,     0, ":*:B::B::::::W::"),
	(0,     0,     0,     '*',     6,     0, ":*:B::B::::::W::"),
	(0,     0,     0,     ':',     4,     0, ":*:B::B::::::W::"),
	(0,     0,     1,     ':',     2,     0, ":*:B::B::::::W::"),
	(0,     0,     1,     'W',     12,     0, ":*:B::B::::::W::"),
	(0,     0,     0,     'B',     15,     0, ":*:B::B:::::WW::"),
	(0,     0,     1,     ':',     11,     0, ":*:B::B:::::WW::"),
	(0,     0,     0,     ':',     10,     0, ":*:B::B:::::WW::"),
	(0,     1,     1,     ':',     1,     0, ":*:B::B:::::WW::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     15,     0, "::::::::::::W:::"),
	(0,     0,     0,     '*',     10,     0, "::::::::::::W::*"),
	(0,     0,     0,     ':',     15,     0, "::::::::::::W::*"),
	(0,     0,     0,     'W',     10,     0, "::::::::::::W::*"),
	(0,     0,     0,     'W',     14,     0, "::::::::::::W::*"),
	(0,     0,     1,     ':',     8,     0, "::::::::::::W::*"),
	(0,     0,     1,     'W',     15,     0, "::::::::::::W::*"),
	(0,     0,     1,     '*',     12,     0, "::::::::::::W::W"),
	(0,     0,     1,     'B',     2,     0, "::::::::::::B::W"),
	(0,     1,     0,     ':',     2,     0, "::B:::::::::B::W"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     2,     0, "::W:::::::::::::"),
	(0,     0,     0,     ':',     4,     0, "::W:::::::::::::"),
	(0,     0,     0,     'W',     6,     0, "::W:::::::::::::"),
	(0,     0,     1,     '*',     0,     0, "::W:::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "*:W:::::::::::::"),
	(0,     0,     0,     '*',     15,     0, "*:W:::::::::::::"),
	(0,     0,     0,     '*',     15,     0, "*:W:::::::::::::"),
	(0,     0,     0,     'B',     9,     0, "*:W:::::::::::::"),
	(0,     0,     0,     'W',     8,     0, "*:W:::::::::::::"),
	(0,     0,     0,     'B',     2,     0, "*:W:::::::::::::"),
	(0,     0,     1,     ':',     8,     0, "*:W:::::::::::::"),
	(0,     1,     0,     'W',     8,     0, "*:W:::::::::::::"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     0, "::W:::::::::::::"),
	(0,     0,     0,     'W',     14,     0, "::W:::::::::::::"),
	(0,     0,     1,     '*',     9,     0, "::W:::::::::::::"),
	(0,     0,     0,     'W',     13,     0, "::W::::::*::::::"),
	(0,     0,     0,     'B',     5,     0, "::W::::::*::::::"),
	(0,     0,     0,     ':',     6,     0, "::W::::::*::::::"),
	(0,     0,     1,     '*',     4,     0, "::W::::::*::::::"),
	(0,     0,     0,     '*',     8,     0, "::W:*::::*::::::"),
	(0,     0,     1,     ':',     5,     0, "::W:*::::*::::::"),
	(0,     0,     1,     'W',     5,     0, "::W:*::::*::::::"),
	(0,     0,     0,     'W',     5,     0, "::W:*W:::*::::::"),
	(0,     0,     1,     ':',     0,     0, "::W:*W:::*::::::"),
	(0,     0,     1,     'B',     8,     0, "::W:*W:::*::::::"),
	(0,     1,     1,     '*',     1,     0, "::W:*W::B*::::::"),
	(0,     0,     0,     'W',     9,     0, ":*::::::::::::::"),
	(0,     0,     0,     'W',     2,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     5,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, ":*:::B::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":*:::B::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":*:::B::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     14,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     3,     0, ":::::B::::::::*:"),
	(0,     0,     1,     'B',     10,     0, ":::B:B::::::::*:"),
	(0,     1,     1,     '*',     11,     0, ":::B:B::::B:::*:"),
	(0,     0,     0,     'B',     2,     0, ":::::::::::*::::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::*::::"),
	(0,     0,     0,     '*',     2,     0, ":::::::::::*::::"),
	(0,     0,     0,     'W',     8,     0, ":::::::::::*::::"),
	(1,     0,     0,     '*',     15,     0, ":::::::::::*::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     14,     0, ":::::W::::::::::"),
	(0,     0,     0,     'B',     15,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     0,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     4,     0, ":::::W:::::::::W"),
	(0,     0,     1,     ':',     0,     0, ":::::W:::::::::W"),
	(0,     0,     0,     '*',     1,     0, ":::::W:::::::::W"),
	(0,     0,     1,     ':',     11,     0, ":::::W:::::::::W"),
	(0,     0,     0,     'W',     11,     0, ":::::W:::::::::W"),
	(0,     0,     1,     'W',     13,     0, ":::::W:::::::::W"),
	(0,     0,     1,     'W',     9,     0, ":::::W:::::::W:W"),
	(0,     0,     1,     '*',     12,     0, ":::::W:::W:::W:W"),
	(0,     0,     1,     ':',     13,     0, ":::::W:::W::*W:W"),
	(0,     1,     1,     ':',     0,     0, ":::::W:::W::*W:W"),
	(0,     0,     0,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     0, ":W::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, ":W::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":W::::::B:::::::"),
	(0,     0,     0,     '*',     10,     0, ":W::::::B:::::::"),
	(0,     0,     0,     '*',     11,     0, ":W::::::B:::::::"),
	(0,     0,     0,     'B',     2,     0, ":W::::::B:::::::"),
	(0,     0,     0,     '*',     1,     0, ":W::::::B:::::::"),
	(0,     0,     0,     'W',     10,     0, ":W::::::B:::::::"),
	(0,     0,     1,     'W',     2,     0, ":W::::::B:::::::"),
	(0,     0,     1,     ':',     9,     0, ":WW:::::B:::::::"),
	(0,     1,     1,     '*',     2,     0, ":WW:::::B:::::::"),
	(0,     0,     0,     ':',     6,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     3,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     13,     0, "::*:::::::::::::"),
	(0,     1,     1,     '*',     13,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     0,     0, ":::::::::::::*::"),
	(0,     0,     1,     ':',     4,     0, ":::::::::::::*::"),
	(0,     0,     1,     '*',     3,     0, ":::::::::::::*::"),
	(0,     0,     1,     ':',     11,     0, ":::*:::::::::*::"),
	(0,     0,     1,     'W',     7,     0, ":::*:::::::::*::"),
	(0,     0,     1,     '*',     6,     0, ":::*:::W:::::*::"),
	(0,     0,     1,     '*',     15,     0, ":::*::*W:::::*::"),
	(0,     0,     1,     'B',     8,     0, ":::*::*W:::::*:*"),
	(0,     0,     1,     'B',     10,     0, ":::*::*WB::::*:*"),
	(0,     0,     0,     ':',     0,     0, ":::*::*WB:B::*:*"),
	(0,     0,     0,     '*',     8,     0, ":::*::*WB:B::*:*"),
	(0,     0,     1,     '*',     13,     0, ":::*::*WB:B::*:*"),
	(0,     0,     0,     ':',     6,     0, ":::*::*WB:B::::*"),
	(0,     0,     0,     'B',     8,     0, ":::*::*WB:B::::*"),
	(0,     0,     0,     ':',     4,     0, ":::*::*WB:B::::*"),
	(0,     0,     0,     ':',     6,     0, ":::*::*WB:B::::*"),
	(0,     0,     1,     '*',     8,     0, ":::*::*WB:B::::*"),
	(0,     1,     1,     '*',     13,     0, ":::*::*WW:B::::*"),
	(0,     0,     1,     'B',     2,     0, ":::::::::::::*::"),
	(0,     0,     1,     ':',     10,     0, "::B::::::::::*::"),
	(0,     0,     0,     'B',     8,     0, "::B::::::::::*::"),
	(0,     0,     0,     'B',     1,     0, "::B::::::::::*::"),
	(0,     0,     0,     'W',     0,     0, "::B::::::::::*::"),
	(0,     0,     1,     ':',     12,     0, "::B::::::::::*::"),
	(0,     0,     0,     'B',     0,     0, "::B::::::::::*::"),
	(0,     0,     1,     'B',     0,     0, "::B::::::::::*::"),
	(0,     1,     1,     ':',     10,     0, "B:B::::::::::*::"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::::::::W:::::"),
	(0,     1,     1,     '*',     0,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     6,     0, "*:::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     5,     0, "*:::::::::::::::"),
	(0,     0,     0,     'B',     2,     0, "*:::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, "*:::::::::::::::"),
	(0,     0,     1,     'W',     10,     0, "*:::::::::::::::"),
	(0,     1,     1,     'B',     9,     0, "*:::::::::W:::::"),
	(0,     0,     1,     ':',     15,     0, ":::::::::B::::::"),
	(0,     0,     1,     '*',     1,     0, ":::::::::B::::::"),
	(0,     0,     0,     ':',     15,     0, ":*:::::::B::::::"),
	(0,     0,     1,     ':',     2,     0, ":*:::::::B::::::"),
	(0,     0,     0,     'B',     3,     0, ":*:::::::B::::::"),
	(0,     0,     1,     'B',     11,     0, ":*:::::::B::::::"),
	(0,     0,     0,     ':',     12,     0, ":*:::::::B:B::::"),
	(0,     0,     0,     '*',     4,     0, ":*:::::::B:B::::"),
	(0,     0,     0,     'B',     7,     0, ":*:::::::B:B::::"),
	(0,     0,     0,     'W',     7,     0, ":*:::::::B:B::::"),
	(0,     0,     1,     '*',     5,     0, ":*:::::::B:B::::"),
	(0,     0,     1,     '*',     3,     0, ":*:::*:::B:B::::"),
	(0,     0,     1,     '*',     0,     0, ":*:*:*:::B:B::::"),
	(0,     0,     0,     'W',     6,     0, "**:*:*:::B:B::::"),
	(0,     0,     1,     '*',     4,     0, "**:*:*:::B:B::::"),
	(0,     0,     0,     'W',     9,     0, "**:***:::B:B::::"),
	(0,     0,     1,     ':',     13,     0, "**:***:::B:B::::"),
	(0,     0,     0,     '*',     8,     0, "**:***:::B:B::::"),
	(0,     0,     1,     'W',     13,     0, "**:***:::B:B::::"),
	(0,     0,     1,     'W',     12,     0, "**:***:::B:B:W::"),
	(0,     0,     0,     ':',     6,     0, "**:***:::B:BWW::"),
	(0,     0,     0,     'B',     7,     0, "**:***:::B:BWW::"),
	(0,     0,     0,     'W',     8,     0, "**:***:::B:BWW::"),
	(0,     0,     1,     'B',     14,     0, "**:***:::B:BWW::"),
	(0,     0,     0,     'W',     14,     0, "**:***:::B:BWWB:"),
	(0,     0,     1,     ':',     15,     0, "**:***:::B:BWWB:"),
	(0,     0,     0,     'W',     10,     0, "**:***:::B:BWWB:"),
	(0,     0,     1,     ':',     2,     0, "**:***:::B:BWWB:"),
	(0,     0,     1,     'B',     13,     0, "**:***:::B:BWWB:"),
	(0,     0,     1,     'B',     1,     0, "**:***:::B:BWBB:"),
	(0,     0,     1,     'W',     5,     0, "*B:***:::B:BWBB:"),
	(0,     0,     0,     'W',     12,     0, "*B:**W:::B:BWBB:"),
	(0,     0,     0,     '*',     8,     0, "*B:**W:::B:BWBB:"),
	(0,     0,     0,     ':',     1,     0, "*B:**W:::B:BWBB:"),
	(0,     1,     0,     '*',     11,     0, "*B:**W:::B:BWBB:"),
	(0,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     14,     0, "::::::W:::::::::"),
	(0,     0,     1,     ':',     0,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     8,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     3,     0, "::::::W:B:::::::"),
	(0,     1,     1,     'B',     8,     0, ":::B::W:B:::::::"),
	(1,     0,     0,     'B',     8,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     0,     0, "B:::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, "B:::::::::::::::"),
	(0,     0,     0,     'W',     3,     0, "B:::::::::::::::"),
	(0,     0,     1,     'W',     10,     0, "B:::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, "B:::::::::W:::::"),
	(0,     0,     0,     '*',     3,     0, "B:::::::::W::::W"),
	(0,     0,     1,     ':',     7,     0, "B:::::::::W::::W"),
	(0,     0,     0,     'W',     12,     0, "B:::::::::W::::W"),
	(0,     1,     1,     '*',     2,     0, "B:::::::::W::::W"),
	(0,     0,     0,     '*',     3,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     6,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     15,     0, "::*:::::::::::::"),
	(0,     1,     0,     'W',     2,     0, "::*:::::::::::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, "::::*:::::::::::"),
	(0,     0,     0,     'W',     12,     0, "*:::*:::::::::::"),
	(0,     0,     0,     '*',     3,     0, "*:::*:::::::::::"),
	(0,     0,     1,     'W',     0,     0, "*:::*:::::::::::"),
	(0,     0,     1,     'W',     9,     0, "W:::*:::::::::::"),
	(0,     0,     1,     '*',     12,     0, "W:::*::::W::::::"),
	(0,     0,     1,     ':',     5,     0, "W:::*::::W::*:::"),
	(0,     0,     0,     'B',     8,     0, "W:::*::::W::*:::"),
	(0,     0,     1,     'B',     5,     0, "W:::*::::W::*:::"),
	(0,     0,     0,     '*',     0,     0, "W:::*B:::W::*:::"),
	(1,     0,     0,     'W',     3,     0, "W:::*B:::W::*:::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::::::::::::B::"),
	(0,     0,     0,     '*',     5,     0, ":::::::::::::B::"),
	(0,     0,     0,     '*',     0,     0, ":::::::::::::B::"),
	(1,     0,     1,     'W',     1,     0, ":::::::::::::B::"),
	(0,     0,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     0, "::::::::::W:::::"),
	(0,     0,     0,     '*',     3,     0, "::::::::::W:::::"),
	(0,     0,     0,     '*',     11,     0, "::::::::::W:::::"),
	(0,     0,     0,     '*',     11,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     15,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     3,     0, "::::::::::W:::::"),
	(1,     1,     0,     '*',     11,     0, "::::::::::W:::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, "::::*:::::::::::"),
	(0,     0,     1,     'W',     10,     0, "::::*:::::::::::"),
	(0,     0,     1,     'W',     4,     0, "::::*:::::W:::::"),
	(0,     0,     1,     ':',     1,     0, "::::W:::::W:::::"),
	(0,     1,     1,     '*',     13,     0, "::::W:::::W:::::"),
	(0,     0,     1,     'W',     2,     0, ":::::::::::::*::"),
	(0,     0,     0,     '*',     15,     0, "::W::::::::::*::"),
	(0,     0,     0,     ':',     12,     0, "::W::::::::::*::"),
	(0,     0,     0,     'W',     11,     0, "::W::::::::::*::"),
	(0,     0,     1,     '*',     15,     0, "::W::::::::::*::"),
	(0,     0,     0,     'B',     2,     0, "::W::::::::::*:*"),
	(0,     1,     1,     ':',     12,     0, "::W::::::::::*:*"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     6,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     2,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     7,     0, "::B:::*:::::::::"),
	(0,     0,     0,     'B',     13,     0, "::B:::**::::::::"),
	(0,     0,     0,     ':',     11,     0, "::B:::**::::::::"),
	(0,     0,     1,     'W',     3,     0, "::B:::**::::::::"),
	(0,     0,     1,     'B',     0,     0, "::BW::**::::::::"),
	(0,     0,     0,     'B',     3,     0, "B:BW::**::::::::"),
	(0,     0,     0,     'B',     13,     0, "B:BW::**::::::::"),
	(0,     0,     0,     'B',     5,     0, "B:BW::**::::::::"),
	(0,     0,     0,     'W',     4,     0, "B:BW::**::::::::"),
	(0,     0,     1,     ':',     10,     0, "B:BW::**::::::::"),
	(0,     0,     1,     ':',     6,     0, "B:BW::**::::::::"),
	(0,     1,     1,     'W',     11,     0, "B:BW::**::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::::::::::W::::"),
	(0,     0,     0,     ':',     11,     0, ":::::::::::W::::"),
	(0,     0,     0,     ':',     11,     0, ":::::::::::W::::"),
	(0,     0,     1,     'B',     11,     0, ":::::::::::W::::"),
	(0,     0,     0,     'W',     7,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     2,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     6,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     13,     0, "::::::B::::B::::"),
	(0,     0,     1,     'B',     11,     0, "::::::B::::B:*::"),
	(0,     0,     1,     'B',     5,     0, "::::::B::::B:*::"),
	(0,     1,     0,     '*',     7,     0, ":::::BB::::B:*::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     12,     0, "B:::::::::::::::"),
	(0,     1,     1,     'W',     13,     0, "B:::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":::::::::::::W::"),
	(0,     0,     0,     ':',     15,     0, ":::::::::::W:W::"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::W:W::"),
	(0,     0,     1,     '*',     15,     0, ":::::::::::W:W::"),
	(0,     0,     1,     'B',     8,     0, ":::::::::::W:W:*"),
	(0,     1,     1,     ':',     2,     0, "::::::::B::W:W:*"),
	(0,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":::::W::::*:::::"),
	(0,     0,     0,     'B',     0,     0, ":::::WW:::*:::::"),
	(0,     0,     1,     ':',     2,     0, ":::::WW:::*:::::"),
	(0,     0,     0,     'B',     15,     0, ":::::WW:::*:::::"),
	(0,     0,     1,     'W',     3,     0, ":::::WW:::*:::::"),
	(0,     0,     0,     'B',     2,     0, ":::W:WW:::*:::::"),
	(0,     0,     1,     'B',     1,     0, ":::W:WW:::*:::::"),
	(1,     0,     1,     'B',     12,     0, ":B:W:WW:::*:::::"),
	(0,     0,     1,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::::::W"),
	(0,     0,     0,     ':',     8,     0, ":::::::::::::::W"),
	(0,     0,     0,     'W',     5,     0, ":::::::::::::::W"),
	(0,     0,     0,     ':',     3,     0, ":::::::::::::::W"),
	(0,     0,     0,     'W',     13,     0, ":::::::::::::::W"),
	(0,     0,     0,     '*',     10,     0, ":::::::::::::::W"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::::::W"),
	(0,     0,     1,     'B',     15,     0, ":::::::::::::::W"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::::::B"),
	(0,     0,     0,     'B',     1,     0, ":::::::::::::::B"),
	(0,     0,     0,     ':',     2,     0, ":::::::::::::::B"),
	(0,     0,     1,     '*',     3,     0, ":::::::::::::::B"),
	(0,     0,     1,     '*',     4,     0, ":::*:::::::::::B"),
	(0,     0,     0,     'B',     3,     0, ":::**::::::::::B"),
	(0,     0,     0,     'B',     2,     0, ":::**::::::::::B"),
	(0,     0,     0,     ':',     9,     0, ":::**::::::::::B"),
	(0,     0,     0,     'B',     3,     0, ":::**::::::::::B"),
	(0,     0,     0,     '*',     1,     0, ":::**::::::::::B"),
	(0,     0,     1,     'W',     4,     0, ":::**::::::::::B"),
	(0,     0,     1,     'B',     14,     0, ":::*W::::::::::B"),
	(0,     0,     0,     ':',     9,     0, ":::*W:::::::::BB"),
	(0,     0,     0,     '*',     15,     0, ":::*W:::::::::BB"),
	(0,     0,     1,     ':',     10,     0, ":::*W:::::::::BB"),
	(0,     1,     1,     '*',     13,     0, ":::*W:::::::::BB"),
	(0,     0,     1,     'W',     1,     0, ":::::::::::::*::"),
	(0,     0,     0,     'W',     2,     0, ":W:::::::::::*::"),
	(0,     0,     1,     ':',     13,     0, ":W:::::::::::*::"),
	(0,     0,     0,     'W',     8,     0, ":W:::::::::::*::"),
	(0,     0,     0,     ':',     2,     0, ":W:::::::::::*::"),
	(0,     1,     0,     '*',     5,     0, ":W:::::::::::*::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     0,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     10,     0, "::::::::B:::::::"),
	(0,     1,     0,     'W',     7,     0, "::::::::B:::::::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "::::::::::::*:::"),
	(0,     0,     1,     ':',     3,     0, "::::W:::::::*:::"),
	(0,     0,     1,     '*',     13,     0, "::::W:::::::*:::"),
	(0,     0,     0,     'W',     4,     0, "::::W:::::::**::"),
	(0,     0,     0,     'B',     11,     0, "::::W:::::::**::"),
	(0,     0,     1,     'W',     11,     0, "::::W:::::::**::"),
	(0,     0,     0,     '*',     4,     0, "::::W::::::W**::"),
	(0,     0,     1,     'W',     4,     0, "::::W::::::W**::"),
	(0,     0,     1,     ':',     0,     0, "::::W::::::W**::"),
	(0,     0,     1,     '*',     0,     0, "::::W::::::W**::"),
	(0,     0,     0,     '*',     14,     0, "*:::W::::::W**::"),
	(0,     0,     0,     'W',     9,     0, "*:::W::::::W**::"),
	(0,     0,     0,     ':',     1,     0, "*:::W::::::W**::"),
	(0,     0,     0,     ':',     15,     0, "*:::W::::::W**::"),
	(0,     0,     1,     'B',     8,     0, "*:::W::::::W**::"),
	(0,     0,     0,     '*',     2,     0, "*:::W:::B::W**::"),
	(0,     0,     0,     'W',     3,     0, "*:::W:::B::W**::"),
	(0,     0,     1,     '*',     15,     0, "*:::W:::B::W**::"),
	(0,     0,     0,     '*',     12,     0, "*:::W:::B::W**:*"),
	(0,     0,     0,     'W',     7,     0, "*:::W:::B::W**:*"),
	(0,     0,     0,     'W',     14,     0, "*:::W:::B::W**:*"),
	(0,     0,     1,     'W',     3,     0, "*:::W:::B::W**:*"),
	(0,     0,     1,     'B',     15,     0, "*::WW:::B::W**:*"),
	(0,     0,     1,     ':',     1,     0, "*::WW:::B::W**:B"),
	(0,     0,     0,     ':',     14,     0, "*::WW:::B::W**:B"),
	(0,     0,     1,     'W',     5,     0, "*::WW:::B::W**:B"),
	(0,     0,     0,     'W',     12,     0, "*::WWW::B::W**:B"),
	(0,     0,     0,     ':',     9,     0, "*::WWW::B::W**:B"),
	(0,     0,     0,     'B',     6,     0, "*::WWW::B::W**:B"),
	(0,     0,     0,     ':',     4,     0, "*::WWW::B::W**:B"),
	(0,     0,     0,     '*',     13,     0, "*::WWW::B::W**:B"),
	(0,     0,     0,     'W',     13,     0, "*::WWW::B::W**:B"),
	(0,     0,     0,     '*',     12,     0, "*::WWW::B::W**:B"),
	(0,     0,     1,     'W',     5,     0, "*::WWW::B::W**:B"),
	(0,     0,     1,     'B',     6,     0, "*::WWW::B::W**:B"),
	(0,     0,     1,     'W',     4,     0, "*::WWWB:B::W**:B"),
	(0,     0,     0,     ':',     4,     0, "*::WWWB:B::W**:B"),
	(0,     1,     0,     ':',     12,     0, "*::WWWB:B::W**:B"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     0, "::::::::::::W:::"),
	(0,     0,     1,     ':',     13,     0, "::::*:::::::W:::"),
	(0,     0,     0,     'W',     14,     0, "::::*:::::::W:::"),
	(0,     0,     1,     'B',     7,     0, "::::*:::::::W:::"),
	(0,     0,     1,     'B',     14,     0, "::::*::B::::W:::"),
	(0,     0,     0,     ':',     0,     0, "::::*::B::::W:B:"),
	(0,     0,     1,     'W',     7,     0, "::::*::B::::W:B:"),
	(0,     0,     1,     ':',     12,     0, "::::*::W::::W:B:"),
	(0,     0,     0,     'B',     5,     0, "::::*::W::::W:B:"),
	(0,     0,     1,     'W',     3,     0, "::::*::W::::W:B:"),
	(0,     0,     1,     'W',     14,     0, ":::W*::W::::W:B:"),
	(0,     0,     1,     ':',     8,     0, ":::W*::W::::W:W:"),
	(0,     1,     0,     'B',     15,     0, ":::W*::W::::W:W:"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     3,     0, "::::*:::::::::::"),
	(0,     0,     0,     'W',     2,     0, "::::*:::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::*:::::::::::"),
	(0,     0,     0,     'W',     15,     0, "::::*:::::::::::"),
	(0,     0,     1,     '*',     10,     0, "::::*:::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::*:::::*:::::"),
	(0,     0,     1,     '*',     6,     0, "::::*:::::*:::::"),
	(0,     0,     1,     'B',     4,     0, "::::*:*:::*:::::"),
	(0,     0,     0,     '*',     12,     0, "::::B:*:::*:::::"),
	(0,     0,     1,     'B',     8,     0, "::::B:*:::*:::::"),
	(0,     0,     0,     '*',     3,     0, "::::B:*:B:*:::::"),
	(0,     0,     0,     '*',     11,     0, "::::B:*:B:*:::::"),
	(1,     0,     0,     '*',     1,     0, "::::B:*:B:*:::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     9,     0, ":::::*::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     15,     0, "::::::::::*:::::"),
	(0,     0,     1,     ':',     4,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     14,     0, ":::::::::::::::B"),
	(0,     0,     0,     ':',     7,     0, ":::::::::::::::B"),
	(0,     1,     1,     '*',     13,     0, ":::::::::::::::B"),
	(0,     1,     1,     'B',     6,     0, ":::::::::::::*::"),
	(0,     0,     0,     'W',     15,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::::B:::::::::"),
	(0,     1,     0,     'W',     12,     0, "::::::B:::::::::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, "::::*:::::::::::"),
	(0,     0,     0,     ':',     15,     0, "::::*:::::::::::"),
	(0,     0,     0,     'W',     7,     0, "::::*:::::::::::"),
	(0,     0,     1,     'W',     4,     0, "::::*:::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     4,     0, "::::W:::::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::B:::::::::::"),
	(0,     0,     1,     '*',     6,     0, "::::B:::::::::::"),
	(0,     0,     1,     'B',     2,     0, "::::B:*:::::::::"),
	(0,     0,     0,     ':',     3,     0, "::B:B:*:::::::::"),
	(0,     0,     1,     '*',     11,     0, "::B:B:*:::::::::"),
	(0,     0,     0,     'B',     7,     0, "::B:B:*::::*::::"),
	(0,     0,     1,     ':',     3,     0, "::B:B:*::::*::::"),
	(0,     0,     0,     ':',     9,     0, "::B:B:*::::*::::"),
	(0,     0,     0,     '*',     6,     0, "::B:B:*::::*::::"),
	(0,     0,     0,     '*',     13,     0, "::B:B:*::::*::::"),
	(0,     1,     0,     ':',     2,     0, "::B:B:*::::*::::"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     8,     0, "::::::W::::W::::"),
	(0,     0,     1,     'B',     11,     0, "::::::W::::W::::"),
	(0,     0,     0,     '*',     0,     0, "::::::W::::B::::"),
	(0,     0,     1,     '*',     5,     0, "::::::W::::B::::"),
	(0,     0,     1,     '*',     15,     0, ":::::*W::::B::::"),
	(0,     0,     0,     'B',     6,     0, ":::::*W::::B:::*"),
	(0,     0,     1,     'W',     6,     0, ":::::*W::::B:::*"),
	(0,     0,     0,     'W',     11,     0, ":::::*W::::B:::*"),
	(0,     0,     0,     'B',     6,     0, ":::::*W::::B:::*"),
	(0,     0,     1,     '*',     9,     0, ":::::*W::::B:::*"),
	(0,     0,     0,     '*',     7,     0, ":::::*W::*:B:::*"),
	(0,     0,     0,     ':',     13,     0, ":::::*W::*:B:::*"),
	(0,     0,     0,     ':',     9,     0, ":::::*W::*:B:::*"),
	(0,     0,     0,     ':',     11,     0, ":::::*W::*:B:::*"),
	(0,     0,     1,     'W',     3,     0, ":::::*W::*:B:::*"),
	(0,     0,     0,     'W',     7,     0, ":::W:*W::*:B:::*"),
	(0,     0,     0,     'W',     3,     0, ":::W:*W::*:B:::*"),
	(0,     0,     1,     ':',     4,     0, ":::W:*W::*:B:::*"),
	(0,     0,     0,     'B',     13,     0, ":::W:*W::*:B:::*"),
	(0,     0,     1,     '*',     12,     0, ":::W:*W::*:B:::*"),
	(0,     0,     0,     '*',     1,     0, ":::W:*W::*:B*::*"),
	(0,     0,     0,     'B',     5,     0, ":::W:*W::*:B*::*"),
	(0,     0,     0,     'W',     15,     0, ":::W:*W::*:B*::*"),
	(0,     0,     0,     'W',     5,     0, ":::W:*W::*:B*::*"),
	(0,     0,     0,     '*',     6,     0, ":::W:*W::*:B*::*"),
	(0,     0,     0,     ':',     15,     0, ":::W:*W::*:B*::*"),
	(0,     0,     1,     'B',     8,     0, ":::W:*W::*:B*::*"),
	(0,     0,     1,     ':',     2,     0, ":::W:*W:B*:B*::*"),
	(0,     1,     0,     ':',     4,     0, ":::W:*W:B*:B*::*"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     13,     0, ":*:::::::::W::::"),
	(0,     1,     1,     'W',     3,     0, ":*:::::::::W::::"),
	(0,     0,     0,     'B',     0,     0, ":::W::::::::::::"),
	(0,     0,     0,     ':',     7,     0, ":::W::::::::::::"),
	(0,     1,     1,     ':',     13,     0, ":::W::::::::::::"),
	(0,     0,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     0,     0, "::::B:::::::::::"),
	(0,     0,     0,     'B',     4,     0, "::::B:::::::::::"),
	(0,     0,     0,     ':',     10,     0, "::::B:::::::::::"),
	(0,     0,     0,     'B',     6,     0, "::::B:::::::::::"),
	(0,     0,     1,     'W',     3,     0, "::::B:::::::::::"),
	(0,     1,     0,     ':',     11,     0, ":::WB:::::::::::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::::::::::::::B"),
	(0,     0,     1,     'W',     4,     0, ":::::::::::::::B"),
	(0,     0,     1,     'B',     2,     0, "::::W::::::::::B"),
	(0,     0,     0,     ':',     5,     0, "::B:W::::::::::B"),
	(0,     0,     0,     'B',     13,     0, "::B:W::::::::::B"),
	(0,     0,     1,     'B',     4,     0, "::B:W::::::::::B"),
	(0,     0,     0,     ':',     8,     0, "::B:B::::::::::B"),
	(0,     0,     0,     'W',     12,     0, "::B:B::::::::::B"),
	(0,     0,     0,     ':',     4,     0, "::B:B::::::::::B"),
	(0,     1,     1,     'B',     9,     0, "::B:B::::::::::B"),
	(0,     0,     0,     '*',     3,     0, ":::::::::B::::::"),
	(0,     0,     0,     ':',     2,     0, ":::::::::B::::::"),
	(0,     0,     1,     'W',     12,     0, ":::::::::B::::::"),
	(0,     0,     1,     'W',     1,     0, ":::::::::B::W:::"),
	(0,     0,     1,     'B',     4,     0, ":W:::::::B::W:::"),
	(0,     0,     1,     'W',     4,     0, ":W::B::::B::W:::"),
	(0,     0,     1,     '*',     4,     0, ":W::W::::B::W:::"),
	(0,     0,     0,     '*',     1,     0, ":W::B::::B::W:::"),
	(0,     0,     0,     'W',     9,     0, ":W::B::::B::W:::"),
	(0,     0,     1,     'W',     2,     0, ":W::B::::B::W:::"),
	(0,     0,     0,     'W',     15,     0, ":WW:B::::B::W:::"),
	(0,     0,     0,     'B',     15,     0, ":WW:B::::B::W:::"),
	(0,     0,     0,     'B',     3,     0, ":WW:B::::B::W:::"),
	(0,     0,     0,     '*',     3,     0, ":WW:B::::B::W:::"),
	(0,     0,     1,     '*',     2,     0, ":WW:B::::B::W:::"),
	(0,     0,     1,     'B',     10,     0, ":WB:B::::B::W:::"),
	(0,     1,     0,     '*',     12,     0, ":WB:B::::BB:W:::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     6,     0, ":::::::::::::W::"),
	(0,     0,     1,     'B',     10,     0, "::::::B:::::::::"),
	(0,     0,     1,     'B',     0,     0, "::::::B:::B:::::"),
	(0,     0,     1,     '*',     10,     0, "B:::::B:::B:::::"),
	(0,     0,     1,     'B',     10,     0, "B:::::B:::W:::::"),
	(0,     0,     1,     '*',     14,     0, "B:::::B:::B:::::"),
	(0,     0,     1,     'W',     10,     0, "B:::::B:::B:::*:"),
	(0,     0,     1,     ':',     3,     0, "B:::::B:::W:::*:"),
	(0,     0,     1,     'W',     0,     0, "B:::::B:::W:::*:"),
	(0,     0,     1,     'W',     12,     0, "W:::::B:::W:::*:"),
	(0,     0,     1,     'W',     15,     0, "W:::::B:::W:W:*:"),
	(0,     0,     1,     '*',     9,     0, "W:::::B:::W:W:*W"),
	(0,     0,     0,     'W',     15,     0, "W:::::B::*W:W:*W"),
	(0,     0,     0,     '*',     7,     0, "W:::::B::*W:W:*W"),
	(0,     0,     1,     ':',     10,     0, "W:::::B::*W:W:*W"),
	(0,     0,     1,     '*',     13,     0, "W:::::B::*W:W:*W"),
	(0,     0,     0,     ':',     0,     0, "W:::::B::*W:W**W"),
	(0,     0,     1,     ':',     3,     0, "W:::::B::*W:W**W"),
	(0,     0,     0,     ':',     10,     0, "W:::::B::*W:W**W"),
	(0,     0,     1,     ':',     1,     0, "W:::::B::*W:W**W"),
	(0,     0,     1,     'W',     11,     0, "W:::::B::*W:W**W"),
	(0,     0,     0,     '*',     7,     0, "W:::::B::*WWW**W"),
	(0,     0,     0,     '*',     8,     0, "W:::::B::*WWW**W"),
	(0,     0,     1,     'W',     4,     0, "W:::::B::*WWW**W"),
	(0,     0,     0,     'W',     5,     0, "W:::W:B::*WWW**W"),
	(0,     0,     0,     ':',     7,     0, "W:::W:B::*WWW**W"),
	(0,     0,     0,     '*',     5,     0, "W:::W:B::*WWW**W"),
	(0,     0,     0,     'W',     12,     0, "W:::W:B::*WWW**W"),
	(0,     0,     1,     'B',     10,     0, "W:::W:B::*WWW**W"),
	(0,     1,     1,     'W',     0,     0, "W:::W:B::*BWW**W"),
	(0,     0,     0,     'W',     13,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     8,     0, "W:::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "W:::::::*:::::::"),
	(0,     0,     0,     'B',     7,     0, "W:::::::*:::::::"),
	(0,     0,     1,     ':',     4,     0, "W:::::::*:::::::"),
	(0,     0,     0,     ':',     3,     0, "W:::::::*:::::::"),
	(0,     0,     0,     'W',     4,     0, "W:::::::*:::::::"),
	(0,     0,     1,     'W',     0,     0, "W:::::::*:::::::"),
	(0,     0,     1,     'B',     12,     0, "W:::::::*:::::::"),
	(0,     0,     1,     'B',     13,     0, "W:::::::*:::B:::"),
	(0,     0,     0,     ':',     5,     0, "W:::::::*:::BB::"),
	(0,     0,     0,     ':',     10,     0, "W:::::::*:::BB::"),
	(0,     0,     1,     'W',     4,     0, "W:::::::*:::BB::"),
	(0,     0,     1,     '*',     3,     0, "W:::W:::*:::BB::"),
	(0,     1,     1,     '*',     13,     0, "W::*W:::*:::BB::"),
	(0,     0,     1,     '*',     10,     0, ":::::::::::::*::"),
	(0,     0,     0,     '*',     13,     0, "::::::::::*::*::"),
	(0,     0,     1,     'B',     2,     0, "::::::::::*::*::"),
	(0,     0,     0,     '*',     0,     0, "::B:::::::*::*::"),
	(0,     0,     1,     'B',     8,     0, "::B:::::::*::*::"),
	(0,     0,     0,     '*',     7,     0, "::B:::::B:*::*::"),
	(0,     0,     0,     'B',     3,     0, "::B:::::B:*::*::"),
	(0,     0,     0,     'B',     5,     0, "::B:::::B:*::*::"),
	(0,     0,     0,     'B',     1,     0, "::B:::::B:*::*::"),
	(0,     0,     1,     'B',     13,     0, "::B:::::B:*::*::"),
	(0,     0,     1,     'W',     0,     0, "::B:::::B:*::B::"),
	(0,     0,     1,     'W',     3,     0, "W:B:::::B:*::B::"),
	(0,     0,     0,     ':',     6,     0, "W:BW::::B:*::B::"),
	(0,     0,     1,     'W',     14,     0, "W:BW::::B:*::B::"),
	(0,     0,     0,     'W',     2,     0, "W:BW::::B:*::BW:"),
	(0,     0,     0,     '*',     0,     0, "W:BW::::B:*::BW:"),
	(0,     0,     1,     '*',     12,     0, "W:BW::::B:*::BW:"),
	(0,     0,     0,     '*',     1,     0, "W:BW::::B:*:*BW:"),
	(0,     0,     0,     ':',     12,     0, "W:BW::::B:*:*BW:"),
	(0,     0,     1,     '*',     2,     0, "W:BW::::B:*:*BW:"),
	(0,     0,     1,     'B',     2,     0, "W:WW::::B:*:*BW:"),
	(0,     0,     0,     'W',     3,     0, "W:BW::::B:*:*BW:"),
	(0,     0,     0,     '*',     8,     0, "W:BW::::B:*:*BW:"),
	(0,     0,     1,     'W',     15,     0, "W:BW::::B:*:*BW:"),
	(0,     0,     1,     'B',     5,     0, "W:BW::::B:*:*BWW"),
	(0,     0,     0,     ':',     10,     0, "W:BW:B::B:*:*BWW"),
	(0,     1,     0,     ':',     9,     0, "W:BW:B::B:*:*BWW"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     0, "::::::::::::*:::"),
	(0,     1,     0,     'B',     10,     0, "::::::::::::*:::"),
	(0,     1,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":::B::::::::::::"),
	(0,     0,     1,     ':',     1,     0, ":::B::::::::::::"),
	(0,     0,     0,     'W',     5,     0, ":::B::::::::::::"),
	(0,     0,     1,     '*',     9,     0, ":::B::::::::::::"),
	(0,     0,     0,     ':',     14,     0, ":::B:::::*::::::"),
	(0,     0,     1,     'B',     1,     0, ":::B:::::*::::::"),
	(0,     0,     1,     ':',     7,     0, ":B:B:::::*::::::"),
	(0,     0,     0,     'B',     7,     0, ":B:B:::::*::::::"),
	(0,     0,     1,     'B',     5,     0, ":B:B:::::*::::::"),
	(0,     0,     0,     'B',     8,     0, ":B:B:B:::*::::::"),
	(0,     1,     1,     '*',     6,     0, ":B:B:B:::*::::::"),
	(0,     0,     0,     '*',     4,     0, "::::::*:::::::::"),
	(0,     0,     1,     'B',     13,     0, "::::::*:::::::::"),
	(0,     0,     1,     'B',     3,     0, "::::::*::::::B::"),
	(0,     0,     0,     '*',     11,     0, ":::B::*::::::B::"),
	(0,     0,     1,     '*',     9,     0, ":::B::*::::::B::"),
	(0,     1,     1,     'W',     1,     0, ":::B::*::*:::B::"),
	(0,     0,     1,     'W',     14,     0, ":W::::::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":W::::::::::::W:"),
	(0,     0,     0,     '*',     5,     0, ":B::::::::::::W:"),
	(0,     0,     0,     ':',     11,     0, ":B::::::::::::W:"),
	(0,     0,     1,     'B',     4,     0, ":B::::::::::::W:"),
	(0,     0,     1,     'B',     13,     0, ":B::B:::::::::W:"),
	(0,     0,     0,     '*',     7,     0, ":B::B::::::::BW:"),
	(0,     0,     0,     ':',     1,     0, ":B::B::::::::BW:"),
	(0,     0,     1,     'B',     7,     0, ":B::B::::::::BW:"),
	(0,     0,     0,     'W',     3,     0, ":B::B::B:::::BW:"),
	(0,     0,     1,     '*',     4,     0, ":B::B::B:::::BW:"),
	(0,     0,     0,     '*',     5,     0, ":B::W::B:::::BW:"),
	(0,     0,     0,     'B',     7,     0, ":B::W::B:::::BW:"),
	(0,     0,     0,     ':',     4,     0, ":B::W::B:::::BW:"),
	(0,     1,     1,     'W',     8,     0, ":B::W::B:::::BW:"),
	(0,     0,     0,     'B',     4,     0, "::::::::W:::::::"),
	(0,     0,     1,     'W',     4,     0, "::::::::W:::::::"),
	(0,     0,     1,     '*',     3,     0, "::::W:::W:::::::"),
	(0,     0,     1,     ':',     9,     0, ":::*W:::W:::::::"),
	(0,     0,     0,     ':',     9,     0, ":::*W:::W:::::::"),
	(0,     0,     0,     'B',     8,     0, ":::*W:::W:::::::"),
	(0,     0,     0,     ':',     15,     0, ":::*W:::W:::::::"),
	(0,     0,     1,     '*',     14,     0, ":::*W:::W:::::::"),
	(0,     0,     1,     '*',     13,     0, ":::*W:::W:::::*:"),
	(0,     0,     1,     ':',     13,     0, ":::*W:::W::::**:"),
	(0,     0,     0,     'B',     15,     0, ":::*W:::W::::**:"),
	(0,     0,     0,     'B',     13,     0, ":::*W:::W::::**:"),
	(0,     0,     0,     'B',     8,     0, ":::*W:::W::::**:"),
	(0,     0,     0,     'W',     14,     0, ":::*W:::W::::**:"),
	(0,     1,     0,     ':',     1,     0, ":::*W:::W::::**:"),
	(0,     0,     0,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::::W:"),
	(0,     0,     0,     'B',     6,     0, "::::::::::::::W:"),
	(0,     0,     0,     '*',     1,     0, "::::::::::::::W:"),
	(0,     0,     0,     '*',     12,     0, "::::::::::::::W:"),
	(0,     1,     1,     '*',     5,     0, "::::::::::::::W:"),
	(0,     0,     1,     'B',     6,     0, ":::::*::::::::::"),
	(0,     1,     1,     'W',     13,     0, ":::::*B:::::::::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::::::W::"),
	(0,     0,     0,     '*',     5,     0, "::::::::*::::W::"),
	(0,     0,     0,     'W',     11,     0, "::::::::*::::W::"),
	(0,     1,     0,     ':',     14,     0, "::::::::*::::W::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     0, ":::::::::::::::B"),
	(0,     0,     1,     ':',     10,     0, "::::::::::::::*B"),
	(0,     0,     0,     'W',     3,     0, "::::::::::::::*B"),
	(0,     0,     1,     ':',     2,     0, "::::::::::::::*B"),
	(0,     0,     0,     '*',     14,     0, "::::::::::::::*B"),
	(0,     0,     0,     'B',     8,     0, "::::::::::::::*B"),
	(0,     0,     1,     'B',     8,     0, "::::::::::::::*B"),
	(0,     0,     1,     'B',     6,     0, "::::::::B:::::*B"),
	(0,     0,     1,     '*',     9,     0, "::::::B:B:::::*B"),
	(0,     0,     1,     'W',     7,     0, "::::::B:B*::::*B"),
	(0,     0,     0,     'B',     12,     0, "::::::BWB*::::*B"),
	(0,     0,     1,     '*',     14,     0, "::::::BWB*::::*B"),
	(0,     0,     1,     '*',     13,     0, "::::::BWB*:::::B"),
	(0,     0,     0,     ':',     13,     0, "::::::BWB*:::*:B"),
	(0,     0,     0,     '*',     1,     0, "::::::BWB*:::*:B"),
	(0,     0,     1,     'B',     13,     0, "::::::BWB*:::*:B"),
	(0,     0,     0,     ':',     5,     0, "::::::BWB*:::B:B"),
	(0,     0,     0,     'W',     6,     0, "::::::BWB*:::B:B"),
	(0,     0,     1,     'B',     2,     0, "::::::BWB*:::B:B"),
	(1,     1,     1,     'W',     12,     0, "::B:::BWB*:::B:B"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, ":::::::::W::::::"),
	(0,     0,     1,     'W',     14,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     5,     0, ":::::::::W::::W:"),
	(0,     0,     0,     '*',     8,     0, ":::::::::W::::W:"),
	(0,     0,     0,     '*',     0,     0, ":::::::::W::::W:"),
	(0,     0,     1,     ':',     14,     0, ":::::::::W::::W:"),
	(0,     0,     0,     '*',     1,     0, ":::::::::W::::W:"),
	(0,     0,     0,     '*',     15,     0, ":::::::::W::::W:"),
	(0,     1,     1,     'W',     11,     0, ":::::::::W::::W:"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::W::::"),
	(0,     0,     1,     '*',     3,     0, ":::::::::::W::::"),
	(0,     0,     0,     '*',     11,     0, ":::*:::::::W::::"),
	(0,     0,     0,     '*',     3,     0, ":::*:::::::W::::"),
	(0,     1,     1,     ':',     0,     0, ":::*:::::::W::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, "::::::B:::::::::"),
	(0,     0,     1,     'B',     9,     0, "::::::B::::B::::"),
	(0,     0,     1,     'W',     10,     0, "::::::B::B:B::::"),
	(0,     0,     1,     ':',     1,     0, "::::::B::BWB::::"),
	(0,     0,     1,     'B',     6,     0, "::::::B::BWB::::"),
	(0,     1,     1,     ':',     11,     0, "::::::B::BWB::::"),
	(0,     1,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     7,     0, "::::::*:::::::::"),
	(0,     1,     0,     'B',     4,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     0, "W:::::::::::::::"),
	(1,     0,     1,     'W',     4,     0, "W::::::::B::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, ":::::::::::*::::"),
	(0,     0,     1,     '*',     11,     0, ":::::::::::*::::"),
	(0,     0,     1,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     12,     0, "::::::::::B:::::"),
	(0,     0,     0,     'W',     7,     0, "::::::::::B:::::"),
	(0,     0,     0,     ':',     2,     0, "::::::::::B:::::"),
	(0,     0,     1,     'B',     14,     0, "::::::::::B:::::"),
	(0,     0,     0,     'W',     7,     0, "::::::::::B:::B:"),
	(0,     0,     1,     '*',     3,     0, "::::::::::B:::B:"),
	(0,     0,     1,     'B',     5,     0, ":::*::::::B:::B:"),
	(0,     0,     1,     ':',     8,     0, ":::*:B::::B:::B:"),
	(0,     0,     0,     'B',     7,     0, ":::*:B::::B:::B:"),
	(0,     0,     0,     '*',     9,     0, ":::*:B::::B:::B:"),
	(0,     0,     0,     ':',     9,     0, ":::*:B::::B:::B:"),
	(0,     0,     1,     'W',     13,     0, ":::*:B::::B:::B:"),
	(0,     0,     0,     'W',     9,     0, ":::*:B::::B::WB:"),
	(0,     0,     1,     '*',     13,     0, ":::*:B::::B::WB:"),
	(0,     0,     1,     'W',     0,     0, ":::*:B::::B::BB:"),
	(0,     0,     0,     '*',     7,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     ':',     7,     0, "W::*:B::::B::BB:"),
	(0,     0,     1,     ':',     4,     0, "W::*:B::::B::BB:"),
	(0,     0,     1,     ':',     11,     0, "W::*:B::::B::BB:"),
	(0,     0,     1,     'B',     13,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     ':',     3,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     '*',     5,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     '*',     0,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     'B',     14,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     ':',     11,     0, "W::*:B::::B::BB:"),
	(1,     0,     0,     'B',     12,     0, "W::*:B::::B::BB:"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     9,     0, "*:::::::::::::::"),
	(0,     1,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, "::::::::W:::::::"),
	(0,     0,     1,     '*',     6,     0, "::::::::W::B::::"),
	(0,     0,     1,     '*',     0,     0, "::::::*:W::B::::"),
	(1,     0,     0,     'B',     3,     0, "*:::::*:W::B::::"),
	(0,     0,     0,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::::*::::::::::"),
	(0,     1,     0,     'W',     8,     0, ":::::*:::::::W::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     7,     0, ":::::::::*::::::"),
	(0,     0,     0,     '*',     15,     0, ":::::::::*::::::"),
	(0,     0,     0,     ':',     8,     0, ":::::::::*::::::"),
	(0,     0,     1,     'B',     11,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     6,     0, ":::::::::*:B::::"),
	(0,     0,     1,     'W',     14,     0, ":::::::::*:B::::"),
	(0,     0,     0,     '*',     7,     0, ":::::::::*:B::W:"),
	(0,     0,     0,     'W',     4,     0, ":::::::::*:B::W:"),
	(0,     0,     1,     '*',     3,     0, ":::::::::*:B::W:"),
	(0,     0,     1,     'W',     7,     0, ":::*:::::*:B::W:"),
	(0,     0,     0,     'B',     11,     0, ":::*:::W:*:B::W:"),
	(0,     0,     0,     '*',     3,     0, ":::*:::W:*:B::W:"),
	(0,     0,     1,     '*',     13,     0, ":::*:::W:*:B::W:"),
	(0,     0,     1,     'B',     10,     0, ":::*:::W:*:B:*W:"),
	(0,     0,     0,     'B',     7,     0, ":::*:::W:*BB:*W:"),
	(0,     0,     0,     '*',     15,     0, ":::*:::W:*BB:*W:"),
	(0,     0,     1,     'W',     8,     0, ":::*:::W:*BB:*W:"),
	(0,     0,     1,     'W',     2,     0, ":::*:::WW*BB:*W:"),
	(0,     0,     0,     '*',     5,     0, "::W*:::WW*BB:*W:"),
	(0,     0,     0,     'B',     5,     0, "::W*:::WW*BB:*W:"),
	(0,     1,     1,     '*',     2,     0, "::W*:::WW*BB:*W:"),
	(0,     0,     1,     ':',     5,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     5,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     13,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     0,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     3,     0, "::*:::::::::::::"),
	(0,     0,     1,     '*',     13,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     10,     0, "::*::::::::::*::"),
	(0,     0,     0,     '*',     15,     0, "::*::::::::::*::"),
	(0,     0,     1,     ':',     6,     0, "::*::::::::::*::"),
	(0,     0,     1,     ':',     0,     0, "::*::::::::::*::"),
	(0,     0,     0,     'B',     2,     0, "::*::::::::::*::"),
	(0,     0,     1,     'B',     14,     0, "::*::::::::::*::"),
	(0,     0,     0,     '*',     10,     0, "::*::::::::::*B:"),
	(0,     0,     1,     'W',     2,     0, "::*::::::::::*B:"),
	(0,     0,     0,     ':',     6,     0, "::W::::::::::*B:"),
	(0,     0,     1,     'B',     15,     0, "::W::::::::::*B:"),
	(0,     0,     1,     ':',     14,     0, "::W::::::::::*BB"),
	(0,     0,     0,     'W',     5,     0, "::W::::::::::*BB"),
	(0,     0,     0,     'B',     12,     0, "::W::::::::::*BB"),
	(0,     0,     0,     ':',     7,     0, "::W::::::::::*BB"),
	(0,     0,     0,     ':',     15,     0, "::W::::::::::*BB"),
	(0,     0,     0,     'B',     9,     0, "::W::::::::::*BB"),
	(0,     0,     0,     'B',     3,     0, "::W::::::::::*BB"),
	(0,     0,     0,     ':',     6,     0, "::W::::::::::*BB"),
	(0,     0,     0,     'W',     11,     0, "::W::::::::::*BB"),
	(0,     0,     1,     '*',     15,     0, "::W::::::::::*BB"),
	(0,     0,     1,     'W',     6,     0, "::W::::::::::*BW"),
	(0,     0,     0,     'B',     13,     0, "::W:::W::::::*BW"),
	(0,     0,     1,     'B',     10,     0, "::W:::W::::::*BW"),
	(0,     0,     0,     ':',     8,     0, "::W:::W:::B::*BW"),
	(0,     0,     1,     ':',     6,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     'B',     7,     0, "::W:::W:::B::*BW"),
	(0,     0,     1,     ':',     0,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     '*',     6,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     'B',     2,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     'B',     0,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     'W',     7,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     ':',     4,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     'B',     15,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     '*',     1,     0, "::W:::W:::B::*BW"),
	(0,     0,     0,     ':',     0,     0, "::W:::W:::B::*BW"),
	(0,     0,     1,     ':',     6,     0, "::W:::W:::B::*BW"),
	(0,     0,     1,     ':',     13,     0, "::W:::W:::B::*BW"),
	(0,     0,     1,     'B',     11,     0, "::W:::W:::B::*BW"),
	(0,     1,     1,     '*',     2,     0, "::W:::W:::BB:*BW"),
	(0,     0,     0,     'B',     4,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     13,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     15,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     3,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     6,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     0,     0, "::*:::B:::::::::"),
	(0,     0,     1,     ':',     6,     0, "::*:::B:::::::::"),
	(0,     1,     1,     'W',     1,     0, "::*:::B:::::::::"),
	(0,     0,     1,     'B',     3,     0, ":W::::::::::::::"),
	(0,     0,     1,     'B',     4,     0, ":W:B::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":W:BB:::::::::::"),
	(0,     0,     0,     '*',     5,     0, ":W:BB:::::::::::"),
	(0,     0,     0,     ':',     12,     0, ":W:BB:::::::::::"),
	(0,     0,     0,     '*',     3,     0, ":W:BB:::::::::::"),
	(0,     0,     1,     'W',     3,     0, ":W:BB:::::::::::"),
	(0,     1,     1,     ':',     14,     0, ":W:WB:::::::::::"),
	(0,     0,     0,     'B',     15,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     1,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     9,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     2,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     7,     0, "::W:::*:::::::::"),
	(0,     0,     1,     '*',     5,     0, "::W:::*:::::::::"),
	(0,     0,     1,     'B',     3,     0, "::W::**:::::::::"),
	(0,     0,     0,     '*',     8,     0, "::WB:**:::::::::"),
	(0,     0,     1,     ':',     10,     0, "::WB:**:::::::::"),
	(0,     0,     0,     ':',     9,     0, "::WB:**:::::::::"),
	(0,     0,     0,     ':',     3,     0, "::WB:**:::::::::"),
	(0,     0,     0,     'W',     14,     0, "::WB:**:::::::::"),
	(0,     0,     0,     ':',     9,     0, "::WB:**:::::::::"),
	(0,     1,     1,     'B',     13,     0, "::WB:**:::::::::"),
	(0,     0,     1,     'W',     3,     0, ":::::::::::::B::"),
	(0,     0,     0,     ':',     8,     0, ":::W:::::::::B::"),
	(0,     0,     1,     'B',     13,     0, ":::W:::::::::B::"),
	(0,     0,     0,     'B',     10,     0, ":::W:::::::::B::"),
	(0,     0,     0,     '*',     10,     0, ":::W:::::::::B::"),
	(0,     0,     0,     'B',     4,     0, ":::W:::::::::B::"),
	(0,     0,     1,     ':',     15,     0, ":::W:::::::::B::"),
	(0,     0,     0,     ':',     10,     0, ":::W:::::::::B::"),
	(0,     0,     0,     'W',     1,     0, ":::W:::::::::B::"),
	(0,     0,     0,     'W',     1,     0, ":::W:::::::::B::"),
	(0,     0,     1,     '*',     2,     0, ":::W:::::::::B::"),
	(0,     1,     1,     'W',     12,     0, "::*W:::::::::B::"),
	(0,     0,     1,     '*',     12,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     6,     0, "::::::::::::B:::"),
	(0,     0,     0,     'B',     8,     0, "::::::::::::B:::"),
	(0,     0,     0,     '*',     15,     0, "::::::::::::B:::"),
	(0,     0,     1,     ':',     0,     0, "::::::::::::B:::"),
	(0,     0,     1,     '*',     3,     0, "::::::::::::B:::"),
	(0,     0,     0,     'B',     4,     0, ":::*::::::::B:::"),
	(0,     0,     1,     'W',     7,     0, ":::*::::::::B:::"),
	(0,     1,     0,     'W',     13,     0, ":::*:::W::::B:::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     12,     0, ":::::::::W::::::"),
	(1,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     15,     0, "::::::::::*:::::"),
	(0,     1,     1,     'W',     4,     0, "::::::::::*::::*"),
	(0,     1,     1,     '*',     2,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     8,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     12,     0, "::*:::::B:::::::"),
	(0,     0,     1,     '*',     8,     0, "::*:::::B:::::::"),
	(0,     0,     1,     'B',     9,     0, "::*:::::W:::::::"),
	(0,     0,     0,     'W',     3,     0, "::*:::::WB::::::"),
	(0,     0,     0,     '*',     13,     0, "::*:::::WB::::::"),
	(0,     0,     1,     ':',     9,     0, "::*:::::WB::::::"),
	(0,     0,     0,     'W',     11,     0, "::*:::::WB::::::"),
	(0,     0,     1,     'B',     1,     0, "::*:::::WB::::::"),
	(0,     1,     1,     'B',     2,     0, ":B*:::::WB::::::"),
	(0,     0,     0,     ':',     5,     0, "::B:::::::::::::"),
	(0,     0,     1,     'W',     7,     0, "::B:::::::::::::"),
	(0,     0,     1,     ':',     5,     0, "::B::::W::::::::"),
	(0,     0,     0,     'B',     13,     0, "::B::::W::::::::"),
	(0,     0,     0,     ':',     0,     0, "::B::::W::::::::"),
	(0,     1,     1,     '*',     2,     0, "::B::::W::::::::"),
	(0,     0,     0,     'B',     15,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     12,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     14,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     5,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::*::W::::::::::"),
	(0,     0,     1,     'W',     11,     0, "::*::W::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::*::W:::::W::::"),
	(0,     1,     0,     'B',     7,     0, "::*::W:::::W::::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     13,     0, "::::B:::::::::B:"),
	(0,     0,     1,     ':',     5,     0, "::::B:::::::::B:"),
	(0,     1,     0,     ':',     11,     0, "::::B:::::::::B:"),
	(0,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     0, ":::::::::::W::::"),
	(0,     0,     0,     'B',     1,     0, ":::::::W:::W::::"),
	(0,     0,     1,     'B',     13,     0, ":::::::W:::W::::"),
	(0,     0,     0,     ':',     7,     0, ":::::::W:::W:B::"),
	(0,     0,     0,     ':',     10,     0, ":::::::W:::W:B::"),
	(0,     0,     1,     ':',     11,     0, ":::::::W:::W:B::"),
	(0,     0,     0,     '*',     1,     0, ":::::::W:::W:B::"),
	(0,     0,     1,     '*',     7,     0, ":::::::W:::W:B::"),
	(0,     0,     0,     '*',     10,     0, ":::::::B:::W:B::"),
	(0,     0,     1,     'W',     0,     0, ":::::::B:::W:B::"),
	(0,     0,     0,     'B',     8,     0, "W::::::B:::W:B::"),
	(0,     0,     0,     'W',     10,     0, "W::::::B:::W:B::"),
	(0,     0,     0,     '*',     11,     0, "W::::::B:::W:B::"),
	(0,     0,     1,     'B',     10,     0, "W::::::B:::W:B::"),
	(0,     0,     0,     'W',     1,     0, "W::::::B::BW:B::"),
	(0,     0,     0,     'B',     4,     0, "W::::::B::BW:B::"),
	(0,     0,     1,     'B',     12,     0, "W::::::B::BW:B::"),
	(0,     1,     1,     'B',     6,     0, "W::::::B::BWBB::"),
	(0,     0,     1,     'B',     9,     0, "::::::B:::::::::"),
	(0,     0,     1,     'B',     4,     0, "::::::B::B::::::"),
	(0,     0,     0,     ':',     15,     0, "::::B:B::B::::::"),
	(0,     0,     1,     'B',     12,     0, "::::B:B::B::::::"),
	(0,     0,     1,     'W',     4,     0, "::::B:B::B::B:::"),
	(0,     0,     0,     'W',     2,     0, "::::W:B::B::B:::"),
	(0,     0,     1,     'W',     1,     0, "::::W:B::B::B:::"),
	(0,     0,     0,     'W',     0,     0, ":W::W:B::B::B:::"),
	(0,     0,     0,     'W',     7,     0, ":W::W:B::B::B:::"),
	(0,     0,     1,     'W',     14,     0, ":W::W:B::B::B:::"),
	(0,     0,     0,     '*',     4,     0, ":W::W:B::B::B:W:"),
	(0,     0,     0,     ':',     7,     0, ":W::W:B::B::B:W:"),
	(0,     1,     0,     ':',     4,     0, ":W::W:B::B::B:W:"),
	(0,     1,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     0, "::::::::::W:::::"),
	(0,     0,     1,     'B',     11,     0, "::::::::::W:::::"),
	(0,     0,     1,     ':',     5,     0, "::::::::::WB::::"),
	(0,     0,     1,     '*',     9,     0, "::::::::::WB::::"),
	(0,     0,     0,     '*',     0,     0, ":::::::::*WB::::"),
	(0,     0,     1,     'W',     11,     0, ":::::::::*WB::::"),
	(0,     0,     0,     ':',     3,     0, ":::::::::*WW::::"),
	(0,     0,     0,     '*',     14,     0, ":::::::::*WW::::"),
	(0,     1,     1,     '*',     7,     0, ":::::::::*WW::::"),
	(0,     0,     1,     ':',     5,     0, ":::::::*::::::::"),
	(0,     1,     0,     ':',     6,     0, ":::::::*::::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, "::::::*:::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     0,     0, "::::::*:::B:::::"),
	(0,     0,     1,     '*',     14,     0, "::::::*:::B:::::"),
	(0,     0,     0,     'B',     12,     0, "::::::*:::B:::*:"),
	(0,     1,     0,     'B',     13,     0, "::::::*:::B:::*:"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, ":::::::::W::::::"),
	(0,     0,     1,     ':',     4,     0, ":::::::::W::::::"),
	(0,     0,     0,     'W',     11,     0, ":::::::::W::::::"),
	(0,     0,     1,     'W',     12,     0, ":::::::::W::::::"),
	(0,     0,     1,     'B',     7,     0, ":::::::::W::W:::"),
	(0,     0,     0,     '*',     6,     0, ":::::::B:W::W:::"),
	(0,     0,     1,     'W',     5,     0, ":::::::B:W::W:::"),
	(0,     0,     0,     'B',     12,     0, ":::::W:B:W::W:::"),
	(0,     0,     1,     ':',     15,     0, ":::::W:B:W::W:::"),
	(0,     0,     0,     '*',     12,     0, ":::::W:B:W::W:::"),
	(0,     0,     0,     'W',     0,     0, ":::::W:B:W::W:::"),
	(0,     0,     1,     'W',     5,     0, ":::::W:B:W::W:::"),
	(0,     0,     1,     'W',     15,     0, ":::::W:B:W::W:::"),
	(0,     0,     0,     'B',     5,     0, ":::::W:B:W::W::W"),
	(0,     0,     1,     ':',     2,     0, ":::::W:B:W::W::W"),
	(0,     0,     0,     ':',     8,     0, ":::::W:B:W::W::W"),
	(0,     0,     1,     'W',     6,     0, ":::::W:B:W::W::W"),
	(0,     0,     1,     ':',     6,     0, ":::::WWB:W::W::W"),
	(0,     0,     1,     'B',     0,     0, ":::::WWB:W::W::W"),
	(0,     0,     0,     ':',     15,     0, "B::::WWB:W::W::W"),
	(0,     0,     1,     '*',     11,     0, "B::::WWB:W::W::W"),
	(0,     0,     0,     ':',     7,     0, "B::::WWB:W:*W::W"),
	(0,     0,     0,     '*',     4,     0, "B::::WWB:W:*W::W"),
	(0,     0,     0,     'W',     10,     0, "B::::WWB:W:*W::W"),
	(0,     0,     1,     '*',     7,     0, "B::::WWB:W:*W::W"),
	(0,     0,     1,     ':',     4,     0, "B::::WWW:W:*W::W"),
	(0,     0,     0,     '*',     8,     0, "B::::WWW:W:*W::W"),
	(0,     0,     0,     'B',     13,     0, "B::::WWW:W:*W::W"),
	(0,     0,     1,     'W',     4,     0, "B::::WWW:W:*W::W"),
	(0,     0,     1,     '*',     12,     0, "B:::WWWW:W:*W::W"),
	(0,     0,     1,     'B',     13,     0, "B:::WWWW:W:*B::W"),
	(0,     0,     1,     'B',     3,     0, "B:::WWWW:W:*BB:W"),
	(0,     0,     1,     ':',     5,     0, "B::BWWWW:W:*BB:W"),
	(0,     0,     0,     'B',     10,     0, "B::BWWWW:W:*BB:W"),
	(0,     1,     1,     ':',     8,     0, "B::BWWWW:W:*BB:W"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     3,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     4,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     5,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     0,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     14,     0, "W:*:::::::::::::"),
	(0,     1,     1,     'W',     15,     0, "W:*:::::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::::::W"),
	(0,     0,     1,     ':',     1,     0, ":::::::::::::::W"),
	(0,     0,     1,     ':',     14,     0, ":::::::::::::::W"),
	(0,     1,     1,     'B',     1,     0, ":::::::::::::::W"),
	(0,     0,     0,     'W',     8,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":B::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":B:::::::::::*::"),
	(0,     0,     1,     'B',     11,     0, ":B:::::::::::*::"),
	(0,     0,     1,     '*',     9,     0, ":B:::::::::B:*::"),
	(0,     0,     1,     'B',     4,     0, ":B:::::::*:B:*::"),
	(0,     0,     1,     'B',     8,     0, ":B::B::::*:B:*::"),
	(0,     0,     0,     '*',     10,     0, ":B::B:::B*:B:*::"),
	(0,     0,     1,     '*',     11,     0, ":B::B:::B*:B:*::"),
	(0,     0,     0,     ':',     14,     0, ":B::B:::B*:W:*::"),
	(0,     0,     1,     'B',     13,     0, ":B::B:::B*:W:*::"),
	(0,     0,     1,     '*',     4,     0, ":B::B:::B*:W:B::"),
	(0,     0,     1,     ':',     6,     0, ":B::W:::B*:W:B::"),
	(0,     0,     0,     'B',     10,     0, ":B::W:::B*:W:B::"),
	(0,     0,     0,     '*',     4,     0, ":B::W:::B*:W:B::"),
	(0,     0,     1,     'W',     11,     0, ":B::W:::B*:W:B::"),
	(0,     0,     0,     ':',     3,     0, ":B::W:::B*:W:B::"),
	(0,     1,     1,     ':',     8,     0, ":B::W:::B*:W:B::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     4,     0, ":::::::::*::::::"),
	(0,     0,     1,     'W',     5,     0, "::::*:::::::::::"),
	(0,     0,     1,     ':',     11,     0, "::::*W::::::::::"),
	(0,     0,     1,     ':',     6,     0, "::::*W::::::::::"),
	(0,     0,     0,     '*',     8,     0, "::::*W::::::::::"),
	(0,     0,     1,     '*',     8,     0, "::::*W::::::::::"),
	(0,     0,     1,     'W',     15,     0, "::::*W::*:::::::"),
	(0,     0,     0,     'W',     8,     0, "::::*W::*::::::W"),
	(0,     0,     1,     '*',     9,     0, "::::*W::*::::::W"),
	(0,     0,     0,     'B',     1,     0, "::::*W::**:::::W"),
	(0,     0,     0,     'W',     2,     0, "::::*W::**:::::W"),
	(0,     0,     0,     'W',     9,     0, "::::*W::**:::::W"),
	(0,     0,     1,     'W',     10,     0, "::::*W::**:::::W"),
	(0,     0,     1,     '*',     8,     0, "::::*W::**W::::W"),
	(0,     0,     1,     'W',     5,     0, "::::*W:::*W::::W"),
	(0,     1,     1,     ':',     6,     0, "::::*W:::*W::::W"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::::::::W:::::::"),
	(0,     0,     1,     '*',     14,     0, "::::::::W:::::::"),
	(0,     0,     0,     '*',     9,     0, "::::::::W:::::*:"),
	(0,     0,     0,     '*',     2,     0, "::::::::W:::::*:"),
	(0,     0,     1,     'W',     6,     0, "::::::::W:::::*:"),
	(0,     0,     1,     'W',     7,     0, "::::::W:W:::::*:"),
	(1,     0,     1,     ':',     8,     0, "::::::WWW:::::*:"),
	(0,     0,     1,     ':',     3,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::::::::W"),
	(0,     1,     1,     'B',     5,     0, "::::::::*::::::W"),
	(0,     0,     1,     '*',     15,     0, ":::::B::::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::::B:::::::::*"),
	(0,     0,     0,     'B',     4,     0, ":::::B:::::::::*"),
	(0,     0,     0,     '*',     12,     0, ":::::B:::::::::*"),
	(0,     0,     1,     'B',     15,     0, ":::::B:::::::::*"),
	(1,     0,     1,     'B',     11,     0, ":::::B:::::::::B"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     0, "::::::W:::::::::"),
	(0,     1,     0,     'B',     1,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, "::::B:::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::::B:::::::::::"),
	(0,     0,     1,     '*',     14,     0, "::::B:::::::::::"),
	(0,     0,     1,     ':',     9,     0, "::::B:::::::::*:"),
	(0,     0,     0,     '*',     7,     0, "::::B:::::::::*:"),
	(0,     0,     0,     '*',     7,     0, "::::B:::::::::*:"),
	(0,     0,     0,     'B',     4,     0, "::::B:::::::::*:"),
	(0,     0,     0,     '*',     10,     0, "::::B:::::::::*:"),
	(0,     0,     0,     '*',     4,     0, "::::B:::::::::*:"),
	(0,     0,     0,     'W',     12,     0, "::::B:::::::::*:"),
	(0,     0,     0,     'W',     8,     0, "::::B:::::::::*:"),
	(0,     0,     1,     'B',     10,     0, "::::B:::::::::*:"),
	(0,     0,     1,     ':',     7,     0, "::::B:::::B:::*:"),
	(0,     0,     0,     ':',     15,     0, "::::B:::::B:::*:"),
	(0,     0,     1,     ':',     14,     0, "::::B:::::B:::*:"),
	(0,     0,     0,     'B',     6,     0, "::::B:::::B:::*:"),
	(0,     0,     0,     'B',     3,     0, "::::B:::::B:::*:"),
	(0,     1,     0,     '*',     8,     0, "::::B:::::B:::*:"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     10,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     4,     0, "::::::::::*:W:::"),
	(0,     0,     0,     ':',     8,     0, "::::*:::::*:W:::"),
	(0,     0,     1,     '*',     0,     0, "::::*:::::*:W:::"),
	(0,     0,     0,     'W',     11,     0, "*:::*:::::*:W:::"),
	(0,     0,     1,     ':',     11,     0, "*:::*:::::*:W:::"),
	(0,     0,     1,     'W',     6,     0, "*:::*:::::*:W:::"),
	(0,     0,     1,     '*',     14,     0, "*:::*:W:::*:W:::"),
	(0,     0,     1,     'B',     8,     0, "*:::*:W:::*:W:*:"),
	(0,     0,     1,     'W',     12,     0, "*:::*:W:B:*:W:*:"),
	(0,     0,     0,     'B',     0,     0, "*:::*:W:B:*:W:*:"),
	(0,     1,     1,     'B',     0,     0, "*:::*:W:B:*:W:*:"),
	(0,     0,     0,     '*',     7,     0, "B:::::::::::::::"),
	(0,     0,     1,     'B',     13,     0, "B:::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "B::::::::::::B::"),
	(0,     0,     0,     '*',     12,     0, "B::::::::::::B::"),
	(0,     0,     1,     'W',     6,     0, "B::::::::::::B::"),
	(0,     0,     1,     'W',     9,     0, "B:::::W::::::B::"),
	(0,     0,     1,     'B',     4,     0, "B:::::W::W:::B::"),
	(0,     0,     1,     ':',     8,     0, "B:::B:W::W:::B::"),
	(0,     0,     0,     'B',     1,     0, "B:::B:W::W:::B::"),
	(0,     0,     0,     ':',     0,     0, "B:::B:W::W:::B::"),
	(0,     1,     1,     ':',     4,     0, "B:::B:W::W:::B::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     5,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     9,     0, ":::::W*:::::::::"),
	(0,     0,     0,     '*',     12,     0, ":::::W*:::::::::"),
	(0,     0,     0,     '*',     2,     0, ":::::W*:::::::::"),
	(0,     0,     1,     ':',     5,     0, ":::::W*:::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::::W*:::::::::"),
	(0,     0,     1,     'B',     12,     0, ":::::W*:::::::::"),
	(0,     0,     1,     ':',     3,     0, ":::::W*:::::B:::"),
	(0,     0,     0,     'B',     3,     0, ":::::W*:::::B:::"),
	(0,     0,     1,     ':',     14,     0, ":::::W*:::::B:::"),
	(0,     0,     0,     ':',     7,     0, ":::::W*:::::B:::"),
	(0,     0,     0,     'W',     0,     0, ":::::W*:::::B:::"),
	(0,     0,     1,     ':',     6,     0, ":::::W*:::::B:::"),
	(0,     0,     0,     ':',     3,     0, ":::::W*:::::B:::"),
	(0,     0,     1,     '*',     7,     0, ":::::W*:::::B:::"),
	(0,     0,     1,     '*',     7,     0, ":::::W**::::B:::"),
	(0,     0,     0,     '*',     6,     0, ":::::W*:::::B:::"),
	(0,     0,     1,     '*',     15,     0, ":::::W*:::::B:::"),
	(0,     0,     1,     'B',     9,     0, ":::::W*:::::B::*"),
	(0,     0,     1,     '*',     9,     0, ":::::W*::B::B::*"),
	(0,     0,     0,     '*',     13,     0, ":::::W*::W::B::*"),
	(0,     0,     0,     'B',     4,     0, ":::::W*::W::B::*"),
	(0,     0,     0,     'B',     15,     0, ":::::W*::W::B::*"),
	(0,     1,     1,     'B',     0,     0, ":::::W*::W::B::*"),
	(0,     0,     1,     'B',     3,     0, "B:::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, "B::B::::::::::::"),
	(0,     0,     1,     'W',     3,     0, "B::B::::::::::::"),
	(0,     0,     0,     'B',     1,     0, "B::W::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "B::W::::::::::::"),
	(0,     0,     1,     ':',     10,     0, "B::W::::::::::::"),
	(0,     0,     0,     ':',     9,     0, "B::W::::::::::::"),
	(0,     0,     1,     '*',     6,     0, "B::W::::::::::::"),
	(0,     0,     1,     'B',     7,     0, "B::W::*:::::::::"),
	(0,     0,     1,     'W',     9,     0, "B::W::*B::::::::"),
	(0,     0,     1,     'W',     15,     0, "B::W::*B:W::::::"),
	(0,     0,     1,     '*',     3,     0, "B::W::*B:W:::::W"),
	(0,     0,     1,     'W',     6,     0, "B::B::*B:W:::::W"),
	(0,     0,     1,     '*',     5,     0, "B::B::WB:W:::::W"),
	(0,     0,     0,     ':',     9,     0, "B::B:*WB:W:::::W"),
	(0,     0,     1,     'W',     1,     0, "B::B:*WB:W:::::W"),
	(0,     0,     1,     '*',     15,     0, "BW:B:*WB:W:::::W"),
	(0,     0,     0,     'B',     8,     0, "BW:B:*WB:W:::::B"),
	(0,     0,     1,     ':',     8,     0, "BW:B:*WB:W:::::B"),
	(0,     0,     0,     '*',     10,     0, "BW:B:*WB:W:::::B"),
	(0,     0,     0,     '*',     11,     0, "BW:B:*WB:W:::::B"),
	(0,     0,     0,     '*',     11,     0, "BW:B:*WB:W:::::B"),
	(0,     0,     0,     'W',     7,     0, "BW:B:*WB:W:::::B"),
	(0,     0,     1,     'W',     4,     0, "BW:B:*WB:W:::::B"),
	(0,     1,     1,     'W',     6,     0, "BW:BW*WB:W:::::B"),
	(0,     0,     1,     ':',     12,     0, "::::::W:::::::::"),
	(0,     0,     0,     '*',     1,     0, "::::::W:::::::::"),
	(0,     0,     0,     '*',     12,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     2,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     2,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     0,     0, "::::::W:::::::::"),
	(0,     1,     1,     '*',     14,     0, "W:::::W:::::::::"),
	(0,     1,     0,     'B',     12,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::::::::::W:::::"),
	(0,     0,     0,     '*',     15,     0, "::::::::::W:::::"),
	(0,     0,     1,     'W',     5,     0, "::::::::::W:::::"),
	(0,     0,     1,     'B',     4,     0, ":::::W::::W:::::"),
	(0,     0,     1,     'W',     6,     0, "::::BW::::W:::::"),
	(0,     0,     1,     ':',     10,     0, "::::BWW:::W:::::"),
	(0,     0,     1,     '*',     14,     0, "::::BWW:::W:::::"),
	(0,     0,     0,     'W',     15,     0, "::::BWW:::W:::*:"),
	(0,     0,     1,     'W',     0,     0, "::::BWW:::W:::*:"),
	(0,     0,     0,     'W',     14,     0, "W:::BWW:::W:::*:"),
	(0,     0,     0,     ':',     3,     0, "W:::BWW:::W:::*:"),
	(0,     0,     1,     'B',     4,     0, "W:::BWW:::W:::*:"),
	(0,     1,     1,     'B',     11,     0, "W:::BWW:::W:::*:"),
	(0,     0,     1,     'W',     5,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     0,     0, ":::::W:::::B::::"),
	(0,     0,     1,     '*',     7,     0, ":::::W:::::B::::"),
	(0,     0,     0,     '*',     2,     0, ":::::W:*:::B::::"),
	(0,     0,     1,     'W',     9,     0, ":::::W:*:::B::::"),
	(0,     0,     0,     'B',     6,     0, ":::::W:*:W:B::::"),
	(0,     0,     0,     'B',     0,     0, ":::::W:*:W:B::::"),
	(0,     0,     1,     'B',     12,     0, ":::::W:*:W:B::::"),
	(0,     1,     0,     '*',     9,     0, ":::::W:*:W:BB:::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     0, ":::::::::::::*::"),
	(0,     0,     0,     'B',     5,     0, "::::::::::W::*::"),
	(0,     0,     1,     ':',     13,     0, "::::::::::W::*::"),
	(0,     0,     0,     'W',     4,     0, "::::::::::W::*::"),
	(1,     0,     0,     '*',     12,     0, "::::::::::W::*::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     0, "::::::*:::::::::"),
	(0,     1,     0,     ':',     1,     0, "::::::*:::W:::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::::::::::B:::::"),
	(0,     0,     1,     'W',     2,     0, "::::::::::B:::::"),
	(0,     0,     1,     '*',     3,     0, "::W:::::::B:::::"),
	(1,     0,     0,     '*',     11,     0, "::W*::::::B:::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     15,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     14,     0, ":::::::::::::::*"),
	(0,     0,     0,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     11,     0, ":::::B::::::::::"),
	(0,     0,     1,     ':',     9,     0, ":::::B::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::::B::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":::::B::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":*:::B::::::::::"),
	(0,     0,     1,     'W',     1,     0, ":*:::B::::::::::"),
	(0,     0,     1,     ':',     4,     0, ":W:::B::::::::::"),
	(0,     1,     0,     'B',     2,     0, ":W:::B::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     0, "::::::::::::W:::"),
	(0,     0,     0,     '*',     1,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     2,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     7,     0, "::W:::::::::W:::"),
	(0,     0,     0,     '*',     3,     0, "::W::::W::::W:::"),
	(0,     0,     1,     ':',     11,     0, "::W::::W::::W:::"),
	(0,     0,     1,     'W',     10,     0, "::W::::W::::W:::"),
	(0,     0,     0,     '*',     4,     0, "::W::::W::W:W:::"),
	(0,     0,     1,     'B',     12,     0, "::W::::W::W:W:::"),
	(0,     0,     0,     ':',     0,     0, "::W::::W::W:B:::"),
	(0,     1,     1,     ':',     5,     0, "::W::::W::W:B:::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     9,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     8,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     14,     0, "::::::::::::W:::"),
	(0,     0,     0,     '*',     2,     0, "::::::::::::W:*:"),
	(0,     0,     0,     '*',     5,     0, "::::::::::::W:*:"),
	(0,     0,     1,     ':',     10,     0, "::::::::::::W:*:"),
	(0,     0,     0,     '*',     5,     0, "::::::::::::W:*:"),
	(0,     0,     0,     '*',     0,     0, "::::::::::::W:*:"),
	(0,     0,     1,     '*',     7,     0, "::::::::::::W:*:"),
	(0,     0,     0,     '*',     11,     0, ":::::::*::::W:*:"),
	(0,     0,     1,     ':',     14,     0, ":::::::*::::W:*:"),
	(0,     0,     0,     'W',     0,     0, ":::::::*::::W:*:"),
	(0,     1,     0,     'W',     0,     0, ":::::::*::::W:*:"),
	(0,     1,     0,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     7,     0, "::::::::::B:W:::"),
	(0,     0,     1,     ':',     10,     0, "::::::::::B:W:::"),
	(0,     0,     1,     '*',     5,     0, "::::::::::B:W:::"),
	(0,     0,     0,     'B',     10,     0, ":::::*::::B:W:::"),
	(0,     0,     0,     ':',     6,     0, ":::::*::::B:W:::"),
	(0,     0,     0,     'B',     3,     0, ":::::*::::B:W:::"),
	(1,     1,     1,     'B',     2,     0, ":::::*::::B:W:::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     6,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     7,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     12,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     10,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     3,     0, "::*:::::::W:::::"),
	(0,     0,     0,     ':',     6,     0, "::*B::::::W:::::"),
	(0,     1,     1,     'W',     7,     0, "::*B::::::W:::::"),
	(1,     0,     1,     ':',     11,     0, ":::::::W::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, "::::::::::W:::::"),
	(0,     0,     1,     '*',     14,     0, "::::::::::W:::::"),
	(0,     1,     0,     ':',     8,     0, "::::::::::W:::*:"),
	(0,     1,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     5,     0, ":*:B::::::::::::"),
	(0,     0,     0,     'W',     14,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     ':',     7,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     'W',     11,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     '*',     11,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     '*',     3,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     '*',     6,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     ':',     2,     0, ":*:B:W::::::::::"),
	(0,     0,     0,     'W',     6,     0, ":*:B:W::::::::::"),
	(0,     1,     1,     'B',     11,     0, ":*:B:W::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     0,     0, ":::::::::::B:W::"),
	(0,     0,     0,     '*',     7,     0, "B::::::::::B:W::"),
	(0,     0,     0,     ':',     1,     0, "B::::::::::B:W::"),
	(0,     0,     1,     ':',     9,     0, "B::::::::::B:W::"),
	(0,     0,     0,     ':',     3,     0, "B::::::::::B:W::"),
	(0,     0,     0,     ':',     2,     0, "B::::::::::B:W::"),
	(0,     0,     1,     'W',     1,     0, "B::::::::::B:W::"),
	(0,     0,     0,     'W',     4,     0, "BW:::::::::B:W::"),
	(0,     0,     1,     'W',     12,     0, "BW:::::::::B:W::"),
	(0,     0,     1,     'B',     6,     0, "BW:::::::::BWW::"),
	(0,     0,     1,     '*',     3,     0, "BW::::B::::BWW::"),
	(0,     0,     1,     'W',     4,     0, "BW:*::B::::BWW::"),
	(0,     0,     1,     'B',     13,     0, "BW:*W:B::::BWW::"),
	(0,     0,     1,     ':',     8,     0, "BW:*W:B::::BWB::"),
	(0,     0,     1,     ':',     9,     0, "BW:*W:B::::BWB::"),
	(0,     0,     1,     'W',     7,     0, "BW:*W:B::::BWB::"),
	(0,     0,     1,     '*',     12,     0, "BW:*W:BW:::BWB::"),
	(0,     0,     0,     '*',     2,     0, "BW:*W:BW:::BBB::"),
	(0,     0,     1,     'B',     14,     0, "BW:*W:BW:::BBB::"),
	(0,     0,     0,     'W',     10,     0, "BW:*W:BW:::BBBB:"),
	(0,     0,     1,     ':',     6,     0, "BW:*W:BW:::BBBB:"),
	(0,     0,     0,     '*',     4,     0, "BW:*W:BW:::BBBB:"),
	(0,     0,     1,     'W',     3,     0, "BW:*W:BW:::BBBB:"),
	(0,     0,     1,     'B',     4,     0, "BW:WW:BW:::BBBB:"),
	(0,     1,     1,     'B',     2,     0, "BW:WB:BW:::BBBB:"),
	(0,     0,     0,     '*',     5,     0, "::B:::::::::::::"),
	(0,     0,     1,     'W',     0,     0, "::B:::::::::::::"),
	(0,     1,     0,     'B',     12,     0, "W:B:::::::::::::"),
	(0,     0,     0,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     15,     0, ":W::::::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":W::::::::::::::"),
	(0,     0,     1,     ':',     1,     0, ":W::::::::::::::"),
	(0,     0,     1,     'B',     2,     0, ":W::::::::::::::"),
	(0,     0,     0,     '*',     2,     0, ":WB:::::::::::::"),
	(0,     0,     1,     'W',     1,     0, ":WB:::::::::::::")
	);
END PACKAGE ex4_data_pak;
