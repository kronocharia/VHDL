
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE WORK.pix_cache_pak.ALL;
USE WORK.pix_tb_pak.ALL;

PACKAGE ex4_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        rst,wen_all,pw: INTEGER;
        pixop:  pixop_tb_t;
        pixnum: INTEGER;
        is_same: INTEGER;
        store: pixop_tb_vec(0 TO 15);
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(
--                 INPUTS              ||           OUTPUTS
--  rst    wen_all  pw   pixop pixnum      is_same   store

	(1,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     0, ":::::::::::::::B"),
	(0,     0,     1,     'B',     3,     0, ":::::::::::::::B"),
	(0,     0,     1,     'B',     9,     0, ":::B:::::::::::B"),
	(0,     1,     1,     'W',     7,     0, ":::B:::::B:::::B"),
	(0,     0,     0,     '*',     11,     0, ":::::::W::::::::"),
	(0,     0,     0,     '*',     11,     0, ":::::::W::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::::::W::::::::"),
	(0,     0,     0,     'B',     3,     0, ":::::::W::::::::"),
	(0,     0,     1,     ':',     10,     0, ":::::::W::::::::"),
	(0,     0,     0,     ':',     10,     0, ":::::::W::::::::"),
	(0,     0,     0,     'B',     12,     0, ":::::::W::::::::"),
	(0,     0,     1,     ':',     7,     0, ":::::::W::::::::"),
	(0,     0,     1,     'W',     4,     0, ":::::::W::::::::"),
	(0,     1,     1,     'B',     1,     0, "::::W::W::::::::"),
	(0,     0,     1,     'B',     3,     0, ":B::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":B:B::::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":B:B::::::::::W:"),
	(0,     0,     1,     'W',     15,     0, ":B:B::::::::::W:"),
	(0,     0,     1,     'B',     13,     0, ":B:B::::::::::WW"),
	(0,     0,     0,     ':',     8,     0, ":B:B:::::::::BWW"),
	(0,     0,     0,     ':',     1,     0, ":B:B:::::::::BWW"),
	(0,     0,     0,     '*',     9,     0, ":B:B:::::::::BWW"),
	(0,     0,     0,     'W',     10,     0, ":B:B:::::::::BWW"),
	(0,     0,     1,     '*',     1,     0, ":B:B:::::::::BWW"),
	(0,     0,     1,     ':',     5,     0, ":W:B:::::::::BWW"),
	(0,     0,     1,     '*',     4,     0, ":W:B:::::::::BWW"),
	(0,     0,     0,     'W',     13,     0, ":W:B*::::::::BWW"),
	(0,     0,     0,     'B',     5,     0, ":W:B*::::::::BWW"),
	(0,     0,     1,     ':',     14,     0, ":W:B*::::::::BWW"),
	(0,     0,     0,     '*',     8,     0, ":W:B*::::::::BWW"),
	(0,     0,     0,     ':',     6,     0, ":W:B*::::::::BWW"),
	(0,     0,     1,     ':',     3,     0, ":W:B*::::::::BWW"),
	(0,     0,     1,     ':',     7,     0, ":W:B*::::::::BWW"),
	(0,     0,     1,     '*',     11,     0, ":W:B*::::::::BWW"),
	(0,     0,     0,     ':',     3,     0, ":W:B*::::::*:BWW"),
	(0,     0,     0,     'B',     3,     0, ":W:B*::::::*:BWW"),
	(0,     0,     0,     ':',     2,     0, ":W:B*::::::*:BWW"),
	(0,     0,     1,     'B',     2,     0, ":W:B*::::::*:BWW"),
	(0,     0,     1,     'B',     10,     0, ":WBB*::::::*:BWW"),
	(0,     0,     1,     '*',     8,     0, ":WBB*:::::B*:BWW"),
	(0,     1,     0,     'B',     0,     0, ":WBB*:::*:B*:BWW"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     0, ":::::::::W::::::"),
	(0,     0,     1,     'W',     13,     0, ":::::::::W::::::"),
	(0,     0,     0,     'W',     4,     0, ":::::::::W:::W::"),
	(0,     1,     0,     'B',     11,     0, ":::::::::W:::W::"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, ":::B::::::::::::"),
	(0,     0,     0,     ':',     5,     0, ":::B::::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::B::::::::::::"),
	(0,     0,     0,     'W',     4,     0, ":::B::::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::B::::::::::::"),
	(0,     0,     1,     'B',     6,     0, ":::B::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::B::B:::::::::"),
	(0,     0,     0,     'W',     12,     0, ":::B::B::::::W::"),
	(0,     1,     0,     'W',     4,     0, ":::B::B::::::W::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":B::::::::::::::"),
	(0,     1,     0,     '*',     13,     0, ":B:::::::::::::W"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "::::::::::::::B:"),
	(0,     0,     1,     'B',     7,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     14,     0, ":::::::B::::::B:"),
	(0,     1,     0,     'W',     11,     0, ":::::::B::::::B:"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     14,     0, "*:::::::::::::::"),
	(0,     1,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     13,     0, "::W:::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::W::::::::::*::"),
	(0,     0,     0,     '*',     0,     0, "::W::::::::::*::"),
	(0,     0,     1,     ':',     2,     0, "::W::::::::::*::"),
	(0,     0,     1,     ':',     7,     0, "::W::::::::::*::"),
	(0,     0,     0,     '*',     7,     0, "::W::::::::::*::"),
	(0,     0,     1,     '*',     12,     0, "::W::::::::::*::"),
	(0,     0,     0,     '*',     2,     0, "::W:::::::::**::"),
	(0,     0,     1,     'W',     6,     0, "::W:::::::::**::"),
	(0,     0,     1,     '*',     0,     0, "::W:::W:::::**::"),
	(0,     0,     1,     'B',     15,     0, "*:W:::W:::::**::"),
	(0,     0,     0,     'B',     3,     0, "*:W:::W:::::**:B"),
	(0,     1,     1,     'W',     14,     0, "*:W:::W:::::**:B"),
	(0,     0,     1,     'B',     2,     0, "::::::::::::::W:"),
	(0,     0,     1,     '*',     11,     0, "::B:::::::::::W:"),
	(0,     0,     0,     '*',     5,     0, "::B::::::::*::W:"),
	(0,     0,     0,     'B',     15,     0, "::B::::::::*::W:"),
	(0,     0,     1,     'W',     10,     0, "::B::::::::*::W:"),
	(0,     0,     1,     'B',     4,     0, "::B:::::::W*::W:"),
	(0,     0,     1,     'B',     2,     0, "::B:B:::::W*::W:"),
	(0,     0,     0,     ':',     10,     0, "::B:B:::::W*::W:"),
	(0,     0,     0,     'B',     9,     0, "::B:B:::::W*::W:"),
	(0,     0,     1,     'B',     4,     0, "::B:B:::::W*::W:"),
	(0,     0,     1,     'W',     1,     0, "::B:B:::::W*::W:"),
	(0,     0,     0,     'B',     15,     0, ":WB:B:::::W*::W:"),
	(0,     0,     0,     ':',     0,     0, ":WB:B:::::W*::W:"),
	(0,     0,     0,     ':',     8,     0, ":WB:B:::::W*::W:"),
	(0,     0,     0,     ':',     5,     0, ":WB:B:::::W*::W:"),
	(0,     0,     1,     '*',     8,     0, ":WB:B:::::W*::W:"),
	(0,     0,     1,     ':',     7,     0, ":WB:B:::*:W*::W:"),
	(0,     0,     0,     ':',     8,     0, ":WB:B:::*:W*::W:"),
	(0,     0,     1,     'B',     8,     0, ":WB:B:::*:W*::W:"),
	(0,     0,     0,     '*',     12,     0, ":WB:B:::B:W*::W:"),
	(0,     0,     1,     '*',     14,     0, ":WB:B:::B:W*::W:"),
	(0,     1,     0,     ':',     6,     0, ":WB:B:::B:W*::B:"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":::::*::::::::::"),
	(0,     1,     1,     ':',     0,     0, ":::::*:::::W::::"),
	(0,     1,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     0, "B:::::::::::::::"),
	(0,     1,     0,     'W',     6,     0, "B:::::::::::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "::B:::::::::::::"),
	(0,     1,     1,     'B',     9,     0, "::B:::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::::::::B::::::"),
	(0,     0,     1,     'B',     3,     0, ":::::::::B:::W::"),
	(0,     0,     1,     'W',     6,     0, ":::B:::::B:::W::"),
	(0,     0,     0,     '*',     7,     0, ":::B::W::B:::W::"),
	(0,     0,     1,     'W',     8,     0, ":::B::W::B:::W::"),
	(0,     0,     0,     'W',     4,     0, ":::B::W:WB:::W::"),
	(0,     0,     0,     ':',     6,     0, ":::B::W:WB:::W::"),
	(0,     0,     0,     'B',     5,     0, ":::B::W:WB:::W::"),
	(0,     0,     0,     'W',     11,     0, ":::B::W:WB:::W::"),
	(0,     0,     0,     '*',     13,     0, ":::B::W:WB:::W::"),
	(0,     0,     0,     '*',     2,     0, ":::B::W:WB:::W::"),
	(0,     0,     1,     '*',     9,     0, ":::B::W:WB:::W::"),
	(0,     0,     1,     'W',     8,     0, ":::B::W:WW:::W::"),
	(0,     0,     1,     'B',     2,     0, ":::B::W:WW:::W::"),
	(0,     0,     1,     ':',     15,     0, "::BB::W:WW:::W::"),
	(0,     1,     0,     '*',     8,     0, "::BB::W:WW:::W::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     3,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     7,     0, ":::W::W:::::::::"),
	(0,     0,     1,     'B',     15,     0, ":::W::WB::::::::"),
	(0,     0,     0,     '*',     15,     0, ":::W::WB:::::::B"),
	(0,     0,     1,     ':',     8,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     'W',     2,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     'B',     5,     0, ":::W::WB:::::::B"),
	(0,     0,     1,     ':',     9,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     '*',     0,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     '*',     5,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     'B',     7,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     'W',     14,     0, ":::W::WB:::::::B"),
	(0,     0,     0,     'B',     7,     0, ":::W::WB:::::::B"),
	(0,     0,     1,     'W',     5,     0, ":::W::WB:::::::B"),
	(0,     1,     0,     '*',     2,     0, ":::W:WWB:::::::B"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     7,     0, ":::::::B::::::::"),
	(0,     0,     1,     '*',     14,     0, ":::::::*::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::::::*::::::*:"),
	(0,     0,     0,     '*',     5,     0, ":::::::*::::::*:"),
	(0,     0,     1,     ':',     13,     0, ":::::::*::::::*:"),
	(0,     0,     1,     ':',     9,     0, ":::::::*::::::*:"),
	(0,     0,     0,     'B',     15,     0, ":::::::*::::::*:"),
	(0,     0,     0,     '*',     4,     0, ":::::::*::::::*:"),
	(0,     0,     0,     ':',     2,     0, ":::::::*::::::*:"),
	(0,     0,     0,     'W',     0,     0, ":::::::*::::::*:"),
	(0,     0,     0,     'B',     0,     0, ":::::::*::::::*:"),
	(0,     0,     0,     '*',     4,     0, ":::::::*::::::*:"),
	(0,     0,     1,     '*',     13,     0, ":::::::*::::::*:"),
	(0,     0,     0,     'W',     1,     0, ":::::::*:::::**:"),
	(0,     0,     1,     ':',     4,     0, ":::::::*:::::**:"),
	(0,     0,     0,     '*',     1,     0, ":::::::*:::::**:"),
	(0,     0,     1,     'W',     13,     0, ":::::::*:::::**:"),
	(0,     0,     0,     ':',     6,     0, ":::::::*:::::W*:"),
	(0,     0,     0,     'W',     10,     0, ":::::::*:::::W*:"),
	(0,     0,     0,     'W',     10,     0, ":::::::*:::::W*:"),
	(0,     0,     0,     'B',     10,     0, ":::::::*:::::W*:"),
	(0,     1,     0,     'B',     11,     0, ":::::::*:::::W*:"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     0, "*:::::::::::::::"),
	(0,     0,     1,     '*',     13,     0, "*B::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, "*B:::::::::::*::"),
	(0,     0,     1,     'B',     4,     0, ":B:::::::::::*::"),
	(0,     0,     1,     '*',     12,     0, ":B::B::::::::*::"),
	(0,     0,     0,     'W',     0,     0, ":B::B:::::::**::"),
	(0,     0,     0,     '*',     0,     0, ":B::B:::::::**::"),
	(0,     0,     0,     'W',     4,     0, ":B::B:::::::**::"),
	(0,     0,     0,     ':',     1,     0, ":B::B:::::::**::"),
	(0,     0,     1,     ':',     3,     0, ":B::B:::::::**::"),
	(0,     1,     1,     '*',     6,     0, ":B::B:::::::**::"),
	(0,     0,     1,     ':',     8,     0, "::::::*:::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     8,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     15,     0, "::::::*:::::::::"),
	(0,     0,     0,     'B',     10,     0, "::::::*::::::::W"),
	(0,     0,     1,     'B',     13,     0, "::::::*::::::::W"),
	(0,     0,     1,     'W',     2,     0, "::::::*::::::B:W"),
	(0,     1,     0,     'W',     5,     0, "::W:::*::::::B:W"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     11,     0, ":::::::::B::::::"),
	(0,     0,     0,     'B',     9,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     10,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     1,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     8,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     0,     0, ":::::::::::B::::"),
	(0,     0,     1,     '*',     6,     0, "B::::::::::B::::"),
	(0,     0,     1,     'B',     14,     0, "B:::::*::::B::::"),
	(0,     0,     0,     'B',     1,     0, "B:::::*::::B::B:"),
	(0,     0,     1,     'W',     11,     0, "B:::::*::::B::B:"),
	(0,     0,     0,     '*',     0,     0, "B:::::*::::W::B:"),
	(0,     0,     0,     'B',     12,     0, "B:::::*::::W::B:"),
	(0,     0,     0,     'W',     13,     0, "B:::::*::::W::B:"),
	(0,     0,     0,     '*',     8,     0, "B:::::*::::W::B:"),
	(0,     0,     0,     '*',     1,     0, "B:::::*::::W::B:"),
	(0,     0,     1,     'W',     13,     0, "B:::::*::::W::B:"),
	(0,     0,     1,     ':',     1,     0, "B:::::*::::W:WB:"),
	(0,     0,     1,     'W',     4,     0, "B:::::*::::W:WB:"),
	(0,     1,     0,     'W',     9,     0, "B:::W:*::::W:WB:"),
	(0,     1,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     2,     0, ":::::::::W::::::"),
	(0,     0,     0,     'B',     8,     0, "::W:::::::::::::"),
	(0,     1,     1,     ':',     1,     0, "::W:::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, ":B::::::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":B::::::B:::::::"),
	(0,     1,     0,     'B',     1,     0, ":B::::::B:::::::"),
	(0,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     2,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     12,     0, "::::::::::::::B:"),
	(0,     0,     0,     ':',     15,     0, "::::::::::::W:B:"),
	(0,     0,     1,     'B',     9,     0, "::::::::::::W:B:"),
	(0,     0,     1,     'B',     9,     0, ":::::::::B::W:B:"),
	(0,     0,     0,     'W',     14,     0, ":::::::::B::W:B:"),
	(0,     0,     0,     '*',     2,     0, ":::::::::B::W:B:"),
	(0,     0,     1,     'W',     11,     0, ":::::::::B::W:B:"),
	(0,     0,     1,     ':',     5,     0, ":::::::::B:WW:B:"),
	(0,     0,     1,     'W',     10,     0, ":::::::::B:WW:B:"),
	(0,     0,     1,     'B',     13,     0, ":::::::::BWWW:B:"),
	(0,     0,     1,     'W',     8,     0, ":::::::::BWWWBB:"),
	(0,     0,     1,     '*',     3,     0, "::::::::WBWWWBB:"),
	(0,     0,     1,     '*',     11,     0, ":::*::::WBWWWBB:"),
	(0,     0,     0,     'W',     4,     0, ":::*::::WBWBWBB:"),
	(0,     1,     0,     'B',     14,     0, ":::*::::WBWBWBB:"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::::::W::::::"),
	(0,     0,     0,     '*',     9,     0, ":::::::::W::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::W::::::"),
	(0,     0,     1,     ':',     8,     0, ":::::::::W::::::"),
	(0,     0,     1,     'B',     12,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::::::W::B:::"),
	(0,     1,     0,     ':',     4,     0, ":::::::::W::B:::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "B:::::::::::W:::"),
	(0,     1,     1,     'B',     11,     0, "B:::::::::::W:::"),
	(0,     0,     1,     'W',     8,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     8,     0, "::::::::W::B::::"),
	(0,     0,     1,     ':',     14,     0, "::::::::W::B::::"),
	(0,     0,     1,     ':',     7,     0, "::::::::W::B::::"),
	(0,     0,     1,     'W',     4,     0, "::::::::W::B::::"),
	(0,     0,     0,     ':',     4,     0, "::::W:::W::B::::"),
	(0,     0,     0,     ':',     6,     0, "::::W:::W::B::::"),
	(0,     0,     0,     'B',     3,     0, "::::W:::W::B::::"),
	(0,     0,     1,     'B',     2,     0, "::::W:::W::B::::"),
	(0,     1,     0,     '*',     11,     0, "::B:W:::W::B::::"),
	(0,     0,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, "::::::::W:::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::::W:::::::"),
	(0,     0,     1,     'W',     15,     0, "::::::::W:::::::"),
	(0,     0,     0,     'W',     6,     0, "::::::::W::::::W"),
	(0,     0,     0,     ':',     11,     0, "::::::::W::::::W"),
	(0,     0,     1,     '*',     13,     0, "::::::::W::::::W"),
	(0,     0,     1,     ':',     2,     0, "::::::::W::::*:W"),
	(0,     0,     0,     'W',     10,     0, "::::::::W::::*:W"),
	(0,     0,     1,     ':',     8,     0, "::::::::W::::*:W"),
	(0,     0,     0,     'W',     11,     0, "::::::::W::::*:W"),
	(0,     0,     0,     ':',     9,     0, "::::::::W::::*:W"),
	(0,     0,     0,     '*',     13,     0, "::::::::W::::*:W"),
	(0,     0,     0,     ':',     0,     0, "::::::::W::::*:W"),
	(0,     0,     0,     '*',     13,     0, "::::::::W::::*:W"),
	(0,     0,     1,     '*',     7,     0, "::::::::W::::*:W"),
	(0,     0,     1,     ':',     9,     0, ":::::::*W::::*:W"),
	(0,     0,     0,     'B',     3,     0, ":::::::*W::::*:W"),
	(0,     0,     0,     ':',     2,     0, ":::::::*W::::*:W"),
	(0,     0,     1,     'B',     6,     0, ":::::::*W::::*:W"),
	(0,     0,     1,     '*',     2,     0, "::::::B*W::::*:W"),
	(0,     0,     1,     '*',     14,     0, "::*:::B*W::::*:W"),
	(0,     0,     0,     'W',     15,     0, "::*:::B*W::::**W"),
	(0,     0,     1,     '*',     5,     0, "::*:::B*W::::**W"),
	(0,     0,     0,     '*',     7,     0, "::*::*B*W::::**W"),
	(0,     0,     1,     'B',     13,     0, "::*::*B*W::::**W"),
	(0,     0,     0,     'B',     8,     0, "::*::*B*W::::B*W"),
	(0,     0,     1,     '*',     13,     0, "::*::*B*W::::B*W"),
	(0,     0,     0,     'W',     2,     0, "::*::*B*W::::W*W"),
	(0,     1,     1,     '*',     3,     0, "::*::*B*W::::W*W"),
	(0,     0,     0,     'B',     1,     0, ":::*::::::::::::"),
	(0,     0,     1,     '*',     6,     0, ":::*::::::::::::"),
	(0,     0,     1,     'W',     1,     0, ":::*::*:::::::::"),
	(0,     0,     1,     'W',     13,     0, ":W:*::*:::::::::"),
	(0,     0,     0,     'W',     14,     0, ":W:*::*::::::W::"),
	(0,     0,     0,     ':',     2,     0, ":W:*::*::::::W::"),
	(0,     0,     0,     ':',     1,     0, ":W:*::*::::::W::"),
	(0,     0,     0,     'W',     15,     0, ":W:*::*::::::W::"),
	(0,     0,     0,     'B',     7,     0, ":W:*::*::::::W::"),
	(0,     0,     1,     '*',     3,     0, ":W:*::*::::::W::"),
	(0,     0,     1,     'B',     2,     0, ":W::::*::::::W::"),
	(0,     1,     0,     ':',     9,     0, ":WB:::*::::::W::"),
	(0,     0,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::::B:::B:::::"),
	(0,     0,     1,     'B',     14,     0, "::::::B:::B:::::"),
	(0,     0,     1,     'W',     2,     0, "::::::B:::B:::B:"),
	(0,     0,     1,     '*',     2,     0, "::W:::B:::B:::B:"),
	(0,     0,     1,     '*',     4,     0, "::B:::B:::B:::B:"),
	(0,     0,     1,     '*',     1,     0, "::B:*:B:::B:::B:"),
	(0,     0,     1,     ':',     10,     0, ":*B:*:B:::B:::B:"),
	(0,     0,     1,     'B',     1,     0, ":*B:*:B:::B:::B:"),
	(0,     0,     1,     'B',     9,     0, ":BB:*:B:::B:::B:"),
	(0,     0,     1,     '*',     7,     0, ":BB:*:B::BB:::B:"),
	(0,     0,     1,     'B',     3,     0, ":BB:*:B*:BB:::B:"),
	(0,     0,     1,     'W',     11,     0, ":BBB*:B*:BB:::B:"),
	(0,     0,     1,     '*',     5,     0, ":BBB*:B*:BBW::B:"),
	(0,     0,     0,     'B',     1,     0, ":BBB**B*:BBW::B:"),
	(0,     1,     1,     'B',     11,     0, ":BBB**B*:BBW::B:"),
	(0,     0,     1,     '*',     7,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     9,     0, ":::::::*:::B::::"),
	(0,     0,     1,     ':',     4,     0, ":::::::*:::B::::"),
	(0,     0,     0,     '*',     11,     0, ":::::::*:::B::::"),
	(0,     0,     0,     ':',     6,     0, ":::::::*:::B::::"),
	(0,     0,     1,     'B',     14,     0, ":::::::*:::B::::"),
	(0,     0,     1,     'B',     3,     0, ":::::::*:::B::B:"),
	(0,     0,     0,     '*',     11,     0, ":::B:::*:::B::B:"),
	(0,     0,     0,     ':',     3,     0, ":::B:::*:::B::B:"),
	(0,     0,     0,     'B',     8,     0, ":::B:::*:::B::B:"),
	(0,     0,     1,     'B',     7,     0, ":::B:::*:::B::B:"),
	(0,     0,     0,     ':',     14,     0, ":::B:::B:::B::B:"),
	(0,     0,     0,     ':',     1,     0, ":::B:::B:::B::B:"),
	(0,     0,     0,     ':',     8,     0, ":::B:::B:::B::B:"),
	(0,     0,     0,     'W',     8,     0, ":::B:::B:::B::B:"),
	(0,     1,     1,     'W',     3,     0, ":::B:::B:::B::B:"),
	(0,     0,     1,     '*',     3,     0, ":::W::::::::::::"),
	(0,     0,     1,     ':',     9,     0, ":::B::::::::::::"),
	(0,     0,     1,     ':',     5,     0, ":::B::::::::::::"),
	(0,     0,     1,     '*',     6,     0, ":::B::::::::::::"),
	(0,     0,     1,     ':',     12,     0, ":::B::*:::::::::"),
	(0,     0,     0,     ':',     3,     0, ":::B::*:::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::B::*:::::::::"),
	(0,     0,     1,     'B',     2,     0, ":::B::*:::::::::"),
	(0,     0,     1,     ':',     10,     0, "::BB::*:::::::::"),
	(0,     0,     0,     'W',     6,     0, "::BB::*:::::::::"),
	(0,     0,     0,     'B',     11,     0, "::BB::*:::::::::"),
	(0,     0,     1,     'B',     5,     0, "::BB::*:::::::::"),
	(0,     0,     1,     'W',     7,     0, "::BB:B*:::::::::"),
	(0,     0,     1,     'W',     4,     0, "::BB:B*W::::::::"),
	(0,     0,     0,     'W',     7,     0, "::BBWB*W::::::::"),
	(0,     0,     1,     ':',     11,     0, "::BBWB*W::::::::"),
	(0,     0,     1,     '*',     12,     0, "::BBWB*W::::::::"),
	(0,     0,     1,     'B',     7,     0, "::BBWB*W::::*:::"),
	(0,     0,     1,     'W',     12,     0, "::BBWB*B::::*:::"),
	(0,     0,     0,     'B',     9,     0, "::BBWB*B::::W:::"),
	(0,     0,     1,     ':',     3,     0, "::BBWB*B::::W:::"),
	(0,     0,     1,     'B',     14,     0, "::BBWB*B::::W:::"),
	(0,     0,     0,     'B',     1,     0, "::BBWB*B::::W:B:"),
	(0,     0,     0,     ':',     0,     0, "::BBWB*B::::W:B:"),
	(0,     1,     0,     'B',     1,     0, "::BBWB*B::::W:B:"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, "::::*:::::::::::"),
	(0,     0,     0,     ':',     12,     0, "::::*:::::::::::"),
	(0,     0,     1,     'B',     3,     0, "::::*:::::::::::"),
	(0,     0,     0,     'B',     10,     0, ":::B*:::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":::B*:::::::::::"),
	(0,     0,     1,     ':',     9,     0, ":::B*::::::W::::"),
	(0,     0,     1,     '*',     9,     0, ":::B*::::::W::::"),
	(0,     0,     0,     ':',     12,     0, ":::B*::::*:W::::"),
	(0,     0,     0,     'W',     11,     0, ":::B*::::*:W::::"),
	(0,     0,     1,     'W',     8,     0, ":::B*::::*:W::::"),
	(0,     0,     1,     ':',     2,     0, ":::B*:::W*:W::::"),
	(0,     0,     0,     '*',     8,     0, ":::B*:::W*:W::::"),
	(0,     0,     0,     'W',     10,     0, ":::B*:::W*:W::::"),
	(0,     0,     0,     '*',     0,     0, ":::B*:::W*:W::::"),
	(0,     0,     0,     ':',     12,     0, ":::B*:::W*:W::::"),
	(0,     0,     1,     '*',     13,     0, ":::B*:::W*:W::::"),
	(0,     0,     0,     ':',     9,     0, ":::B*:::W*:W:*::"),
	(0,     0,     0,     ':',     8,     0, ":::B*:::W*:W:*::"),
	(0,     0,     1,     'W',     13,     0, ":::B*:::W*:W:*::"),
	(0,     0,     1,     'W',     5,     0, ":::B*:::W*:W:W::"),
	(0,     0,     1,     'W',     12,     0, ":::B*W::W*:W:W::"),
	(0,     0,     0,     '*',     11,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     'B',     0,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     '*',     5,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     'B',     9,     0, ":::B*W::W*:WWW::"),
	(0,     0,     1,     'W',     13,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     'W',     10,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     'W',     0,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     '*',     1,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     'W',     2,     0, ":::B*W::W*:WWW::"),
	(0,     0,     1,     ':',     5,     0, ":::B*W::W*:WWW::"),
	(0,     0,     1,     '*',     3,     0, ":::B*W::W*:WWW::"),
	(0,     0,     0,     'B',     13,     0, ":::W*W::W*:WWW::"),
	(0,     0,     0,     ':',     6,     0, ":::W*W::W*:WWW::"),
	(0,     0,     0,     ':',     2,     0, ":::W*W::W*:WWW::"),
	(0,     0,     0,     ':',     8,     0, ":::W*W::W*:WWW::"),
	(0,     0,     0,     'W',     1,     0, ":::W*W::W*:WWW::"),
	(0,     0,     1,     '*',     4,     0, ":::W*W::W*:WWW::"),
	(0,     1,     0,     'W',     15,     0, ":::W:W::W*:WWW::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     12,     0, ":::::B::::::::::"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     13,     0, "::::::::::B:::B:"),
	(0,     1,     0,     '*',     13,     0, "::::::::::B:::B:"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     4,     0, ":::::W::::::::::"),
	(0,     0,     0,     'B',     7,     0, ":::::W::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     7,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     7,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::::W::::::::::"),
	(0,     0,     1,     'W',     5,     0, ":::::W:::::::::W"),
	(0,     0,     0,     'W',     5,     0, ":::::W:::::::::W"),
	(0,     0,     1,     'W',     2,     0, ":::::W:::::::::W"),
	(0,     0,     1,     ':',     5,     0, "::W::W:::::::::W"),
	(0,     0,     1,     ':',     5,     0, "::W::W:::::::::W"),
	(0,     0,     0,     ':',     10,     0, "::W::W:::::::::W"),
	(0,     1,     1,     '*',     2,     0, "::W::W:::::::::W"),
	(0,     0,     0,     'B',     15,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     9,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     15,     0, "::*::::::W::::::"),
	(0,     0,     0,     'W',     7,     0, "::*::::::W:::::W"),
	(0,     0,     0,     'B',     1,     0, "::*::::::W:::::W"),
	(0,     0,     0,     'B',     14,     0, "::*::::::W:::::W"),
	(0,     0,     1,     ':',     8,     0, "::*::::::W:::::W"),
	(0,     0,     1,     '*',     9,     0, "::*::::::W:::::W"),
	(0,     1,     1,     ':',     10,     0, "::*::::::B:::::W"),
	(0,     0,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, ":::::::W::::::::"),
	(0,     0,     1,     ':',     3,     0, "*::::::W::::::::"),
	(0,     0,     1,     'B',     6,     0, "*::::::W::::::::"),
	(0,     0,     0,     ':',     6,     0, "*:::::BW::::::::"),
	(0,     0,     0,     ':',     10,     0, "*:::::BW::::::::"),
	(0,     0,     0,     ':',     7,     0, "*:::::BW::::::::"),
	(0,     0,     1,     ':',     3,     0, "*:::::BW::::::::"),
	(0,     0,     0,     ':',     7,     0, "*:::::BW::::::::"),
	(0,     0,     0,     'W',     7,     0, "*:::::BW::::::::"),
	(0,     0,     1,     '*',     15,     0, "*:::::BW::::::::"),
	(0,     0,     0,     'W',     7,     0, "*:::::BW:::::::*"),
	(0,     0,     0,     'B',     13,     0, "*:::::BW:::::::*"),
	(0,     0,     1,     'B',     0,     0, "*:::::BW:::::::*"),
	(0,     0,     1,     'W',     1,     0, "B:::::BW:::::::*"),
	(0,     1,     1,     'W',     13,     0, "BW::::BW:::::::*"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::::W::"),
	(0,     0,     1,     'B',     2,     0, ":::::::::::::W::"),
	(0,     0,     0,     'W',     3,     0, "::B::::::::::W::"),
	(0,     0,     1,     ':',     0,     0, "::B::::::::::W::"),
	(0,     0,     0,     'B',     13,     0, "::B::::::::::W::"),
	(0,     0,     0,     'B',     15,     0, "::B::::::::::W::"),
	(0,     0,     1,     'W',     1,     0, "::B::::::::::W::"),
	(0,     0,     0,     '*',     7,     0, ":WB::::::::::W::"),
	(0,     0,     0,     '*',     8,     0, ":WB::::::::::W::"),
	(0,     1,     1,     'W',     3,     0, ":WB::::::::::W::"),
	(0,     0,     0,     '*',     15,     0, ":::W::::::::::::"),
	(0,     0,     1,     '*',     11,     0, ":::W::::::::::::"),
	(0,     0,     1,     'W',     8,     0, ":::W:::::::*::::"),
	(0,     0,     0,     ':',     12,     0, ":::W::::W::*::::"),
	(0,     1,     1,     'W',     12,     0, ":::W::::W::*::::"),
	(0,     0,     1,     ':',     15,     0, "::::::::::::W:::"),
	(0,     0,     0,     '*',     10,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     7,     0, "::::::::::::W:::"),
	(0,     0,     1,     ':',     3,     0, "::::::::::::W:::"),
	(0,     0,     0,     'W',     10,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     7,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     9,     0, ":::::::*::::W:::"),
	(0,     0,     1,     'W',     6,     0, ":::::::*::::W:::"),
	(0,     0,     0,     'B',     14,     0, "::::::W*::::W:::"),
	(0,     1,     1,     'B',     11,     0, "::::::W*::::W:::"),
	(0,     0,     1,     'W',     7,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     7,     0, ":::::::W:::B::::"),
	(0,     0,     1,     'W',     11,     0, ":::::::B:::B::::"),
	(0,     0,     1,     '*',     14,     0, ":::::::B:::W::::"),
	(0,     0,     0,     'W',     8,     0, ":::::::B:::W::*:"),
	(0,     0,     0,     ':',     0,     0, ":::::::B:::W::*:"),
	(0,     1,     0,     'W',     7,     0, ":::::::B:::W::*:"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::::::B::"),
	(0,     1,     1,     'W',     13,     0, "::::::::*::::B::"),
	(0,     0,     0,     'B',     5,     0, ":::::::::::::W::"),
	(0,     0,     0,     ':',     2,     0, ":::::::::::::W::"),
	(0,     0,     0,     'W',     3,     0, ":::::::::::::W::"),
	(0,     0,     1,     'W',     12,     0, ":::::::::::::W::"),
	(0,     0,     1,     'B',     13,     0, "::::::::::::WW::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::::WB::"),
	(0,     0,     1,     'W',     2,     0, "::::::::::::WB::"),
	(0,     1,     1,     '*',     5,     0, "::W:::::::::WB::"),
	(0,     0,     0,     'W',     13,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":::::*::::::::::"),
	(0,     0,     1,     'B',     8,     0, ":::::*::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::*::B:::::::"),
	(0,     0,     1,     '*',     10,     0, ":::::*::B:::::::"),
	(0,     1,     1,     'B',     13,     0, ":::::*::B:*:::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::::B::"),
	(0,     0,     1,     'B',     13,     0, ":::::::::::::B::"),
	(0,     0,     1,     'B',     14,     0, ":::::::::::::B::"),
	(0,     0,     0,     'W',     3,     0, ":::::::::::::BB:"),
	(0,     0,     1,     '*',     14,     0, ":::::::::::::BB:"),
	(0,     0,     0,     'W',     2,     0, ":::::::::::::BW:"),
	(0,     0,     1,     'B',     13,     0, ":::::::::::::BW:"),
	(0,     0,     0,     '*',     0,     0, ":::::::::::::BW:"),
	(0,     0,     1,     'B',     2,     0, ":::::::::::::BW:"),
	(0,     0,     1,     'B',     7,     0, "::B::::::::::BW:"),
	(0,     1,     1,     '*',     1,     0, "::B::::B:::::BW:"),
	(0,     0,     0,     'W',     5,     0, ":*::::::::::::::"),
	(0,     0,     1,     '*',     4,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     15,     0, ":*::*:::::::::::"),
	(0,     0,     0,     '*',     0,     0, ":*::*:::::::::::"),
	(0,     1,     1,     ':',     15,     0, ":*::*:::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::*:::::::::::"),
	(0,     0,     0,     '*',     3,     0, "::*:*:::::::::::"),
	(0,     0,     0,     'W',     14,     0, "::*:*:::::::::::"),
	(0,     0,     1,     'B',     3,     0, "::*:*:::::::::::"),
	(0,     0,     0,     'W',     10,     0, "::*B*:::::::::::"),
	(0,     1,     1,     'W',     3,     0, "::*B*:::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":::W::::::::::::"),
	(0,     0,     0,     '*',     0,     0, ":*:W::::::::::::"),
	(0,     0,     1,     '*',     9,     0, ":*:W::::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":*:W:::::*::::::"),
	(0,     0,     0,     'B',     8,     0, ":*:W:::::*::::::"),
	(0,     0,     1,     ':',     10,     0, ":*:W:::::*::::::"),
	(0,     0,     0,     'W',     11,     0, ":*:W:::::*::::::"),
	(0,     0,     0,     '*',     0,     0, ":*:W:::::*::::::"),
	(0,     0,     1,     'B',     5,     0, ":*:W:::::*::::::"),
	(0,     0,     1,     '*',     10,     0, ":*:W:B:::*::::::"),
	(0,     0,     1,     'W',     8,     0, ":*:W:B:::**:::::"),
	(0,     0,     0,     '*',     1,     0, ":*:W:B::W**:::::"),
	(0,     0,     0,     'W',     13,     0, ":*:W:B::W**:::::"),
	(0,     0,     0,     'B',     15,     0, ":*:W:B::W**:::::"),
	(0,     0,     1,     '*',     11,     0, ":*:W:B::W**:::::"),
	(0,     0,     1,     '*',     11,     0, ":*:W:B::W***::::"),
	(0,     0,     1,     'W',     8,     0, ":*:W:B::W**:::::"),
	(0,     0,     0,     'B',     7,     0, ":*:W:B::W**:::::"),
	(0,     0,     1,     '*',     11,     0, ":*:W:B::W**:::::"),
	(0,     0,     0,     'W',     13,     0, ":*:W:B::W***::::"),
	(0,     1,     0,     'W',     5,     0, ":*:W:B::W***::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":::::B::::::::::"),
	(0,     0,     1,     ':',     13,     0, ":::::B::::::*:::"),
	(0,     0,     1,     ':',     5,     0, ":::::B::::::*:::"),
	(0,     0,     1,     '*',     1,     0, ":::::B::::::*:::"),
	(0,     0,     1,     ':',     6,     0, ":*:::B::::::*:::"),
	(0,     0,     1,     'B',     14,     0, ":*:::B::::::*:::"),
	(0,     0,     1,     '*',     15,     0, ":*:::B::::::*:B:"),
	(0,     0,     1,     'W',     1,     0, ":*:::B::::::*:B*"),
	(0,     0,     1,     'B',     2,     0, ":W:::B::::::*:B*"),
	(0,     0,     0,     '*',     5,     0, ":WB::B::::::*:B*"),
	(0,     0,     1,     ':',     8,     0, ":WB::B::::::*:B*"),
	(0,     0,     0,     'W',     0,     0, ":WB::B::::::*:B*"),
	(0,     0,     1,     'W',     13,     0, ":WB::B::::::*:B*"),
	(0,     0,     0,     '*',     4,     0, ":WB::B::::::*WB*"),
	(0,     0,     1,     'W',     1,     0, ":WB::B::::::*WB*"),
	(0,     0,     1,     '*',     8,     0, ":WB::B::::::*WB*"),
	(0,     0,     0,     'W',     15,     0, ":WB::B::*:::*WB*"),
	(0,     0,     0,     '*',     4,     0, ":WB::B::*:::*WB*"),
	(0,     0,     1,     'B',     13,     0, ":WB::B::*:::*WB*"),
	(0,     0,     0,     ':',     4,     0, ":WB::B::*:::*BB*"),
	(0,     0,     0,     'W',     13,     0, ":WB::B::*:::*BB*"),
	(0,     0,     1,     'W',     14,     0, ":WB::B::*:::*BB*"),
	(0,     0,     1,     'W',     0,     0, ":WB::B::*:::*BW*"),
	(0,     0,     1,     ':',     6,     0, "WWB::B::*:::*BW*"),
	(0,     0,     0,     ':',     10,     0, "WWB::B::*:::*BW*"),
	(0,     1,     0,     'W',     13,     0, "WWB::B::*:::*BW*"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::::::::::::*:"),
	(0,     0,     1,     'W',     3,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     10,     0, ":::W::::::::::*:"),
	(0,     0,     0,     ':',     0,     0, ":::W::::::::::*:"),
	(0,     0,     1,     ':',     13,     0, ":::W::::::::::*:"),
	(0,     0,     0,     'W',     11,     0, ":::W::::::::::*:"),
	(0,     0,     0,     'W',     4,     0, ":::W::::::::::*:"),
	(0,     0,     0,     'B',     12,     0, ":::W::::::::::*:"),
	(0,     0,     0,     'W',     5,     0, ":::W::::::::::*:"),
	(0,     0,     1,     '*',     14,     0, ":::W::::::::::*:"),
	(0,     0,     0,     'B',     4,     0, ":::W::::::::::::"),
	(0,     0,     1,     'B',     10,     0, ":::W::::::::::::"),
	(0,     0,     1,     ':',     5,     0, ":::W::::::B:::::"),
	(0,     0,     1,     ':',     2,     0, ":::W::::::B:::::"),
	(0,     0,     1,     '*',     2,     0, ":::W::::::B:::::"),
	(0,     0,     0,     'B',     13,     0, "::*W::::::B:::::"),
	(0,     0,     1,     '*',     9,     0, "::*W::::::B:::::"),
	(0,     1,     1,     'W',     9,     0, "::*W:::::*B:::::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::W::::::"),
	(0,     0,     1,     'B',     6,     0, "::::::::*W::::::"),
	(0,     0,     1,     'B',     2,     0, "::::::B:*W::::::"),
	(0,     0,     0,     'B',     8,     0, "::B:::B:*W::::::"),
	(0,     0,     0,     'B',     3,     0, "::B:::B:*W::::::"),
	(0,     0,     1,     'W',     1,     0, "::B:::B:*W::::::"),
	(0,     0,     1,     ':',     11,     0, ":WB:::B:*W::::::"),
	(0,     0,     1,     'W',     4,     0, ":WB:::B:*W::::::"),
	(0,     0,     1,     '*',     4,     0, ":WB:W:B:*W::::::"),
	(0,     0,     1,     ':',     15,     0, ":WB:B:B:*W::::::"),
	(0,     0,     1,     'W',     11,     0, ":WB:B:B:*W::::::"),
	(0,     0,     1,     'B',     0,     0, ":WB:B:B:*W:W::::"),
	(0,     0,     0,     'W',     9,     0, "BWB:B:B:*W:W::::"),
	(0,     0,     0,     'B',     2,     0, "BWB:B:B:*W:W::::"),
	(0,     0,     1,     ':',     11,     0, "BWB:B:B:*W:W::::"),
	(0,     0,     1,     'W',     7,     0, "BWB:B:B:*W:W::::"),
	(0,     0,     1,     'B',     15,     0, "BWB:B:BW*W:W::::"),
	(0,     1,     1,     ':',     15,     0, "BWB:B:BW*W:W:::B"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     1,     0, ":*::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     7,     0, "::::::::::*:::::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":*::::::::::::::"),
	(0,     0,     0,     ':',     13,     0, ":*::::::::::::::"),
	(0,     0,     1,     '*',     1,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     8,     0, "::::::::::::*:::"),
	(0,     1,     0,     ':',     6,     0, "::::::::W:::*:::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::::::*::::::::"),
	(0,     0,     1,     'B',     4,     0, ":::::::*::::::::"),
	(0,     0,     1,     '*',     0,     0, "::::B::*::::::::"),
	(0,     0,     0,     ':',     13,     0, "*:::B::*::::::::"),
	(0,     0,     1,     'W',     15,     0, "*:::B::*::::::::"),
	(0,     0,     0,     '*',     12,     0, "*:::B::*:::::::W"),
	(0,     0,     1,     '*',     9,     0, "*:::B::*:::::::W"),
	(0,     0,     1,     'W',     13,     0, "*:::B::*:*:::::W"),
	(0,     0,     1,     ':',     12,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     ':',     11,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     'B',     12,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     'W',     9,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     '*',     14,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     ':',     9,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     'B',     13,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     'B',     1,     0, "*:::B::*:*:::W:W"),
	(0,     0,     1,     'W',     5,     0, "*:::B::*:*:::W:W"),
	(0,     0,     0,     '*',     13,     0, "*:::BW:*:*:::W:W"),
	(0,     0,     1,     '*',     15,     0, "*:::BW:*:*:::W:W"),
	(0,     0,     0,     '*',     5,     0, "*:::BW:*:*:::W:B"),
	(0,     0,     1,     ':',     15,     0, "*:::BW:*:*:::W:B"),
	(0,     0,     0,     ':',     5,     0, "*:::BW:*:*:::W:B"),
	(0,     0,     1,     '*',     4,     0, "*:::BW:*:*:::W:B"),
	(0,     0,     1,     'W',     8,     0, "*:::WW:*:*:::W:B"),
	(0,     0,     0,     'B',     14,     0, "*:::WW:*W*:::W:B"),
	(0,     0,     1,     'B',     11,     0, "*:::WW:*W*:::W:B"),
	(0,     0,     0,     '*',     12,     0, "*:::WW:*W*:B:W:B"),
	(0,     1,     1,     '*',     0,     0, "*:::WW:*W*:B:W:B"),
	(0,     0,     1,     'B',     12,     0, "*:::::::::::::::"),
	(0,     0,     1,     '*',     1,     0, "*:::::::::::B:::"),
	(0,     0,     1,     'B',     2,     0, "**::::::::::B:::"),
	(0,     0,     0,     'W',     11,     0, "**B:::::::::B:::"),
	(0,     0,     1,     'W',     0,     0, "**B:::::::::B:::"),
	(0,     0,     1,     'B',     3,     0, "W*B:::::::::B:::"),
	(0,     0,     0,     '*',     14,     0, "W*BB::::::::B:::"),
	(0,     0,     1,     '*',     3,     0, "W*BB::::::::B:::"),
	(0,     1,     1,     '*',     9,     0, "W*BW::::::::B:::"),
	(0,     0,     1,     ':',     6,     0, ":::::::::*::::::"),
	(0,     1,     0,     'W',     3,     0, ":::::::::*::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "::*:::::::::::::"),
	(0,     1,     0,     ':',     4,     0, "::*:W:::::::::::"),
	(0,     0,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     11,     0, "::::::::::::::W:"),
	(0,     0,     0,     'B',     15,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     0,     0, ":::::::::::B::::"),
	(0,     0,     0,     '*',     8,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     3,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     0,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     3,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     3,     0, ":::::::::::B::::"),
	(0,     1,     1,     '*',     2,     0, ":::::::::::B::::"),
	(0,     0,     1,     'W',     9,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     7,     0, "::*::::::W::::::"),
	(0,     1,     1,     'W',     15,     0, "::*::::::W::::::"),
	(0,     0,     1,     '*',     14,     0, ":::::::::::::::W"),
	(0,     0,     1,     'W',     9,     0, "::::::::::::::*W"),
	(0,     0,     0,     'W',     11,     0, ":::::::::W::::*W"),
	(0,     0,     0,     ':',     7,     0, ":::::::::W::::*W"),
	(0,     0,     1,     ':',     6,     0, ":::::::::W::::*W"),
	(0,     1,     0,     '*',     7,     0, ":::::::::W::::*W"),
	(0,     0,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::*:::::::::::W:"),
	(0,     0,     1,     'B',     2,     0, "::*:::::::::::W:"),
	(0,     0,     1,     ':',     5,     0, "::B:::::::::::W:"),
	(0,     0,     0,     'B',     0,     0, "::B:::::::::::W:"),
	(0,     0,     0,     'B',     6,     0, "::B:::::::::::W:"),
	(0,     0,     0,     'B',     2,     0, "::B:::::::::::W:"),
	(0,     0,     1,     'W',     12,     0, "::B:::::::::::W:"),
	(0,     0,     1,     ':',     15,     0, "::B:::::::::W:W:"),
	(0,     0,     1,     'B',     8,     0, "::B:::::::::W:W:"),
	(0,     0,     0,     'B',     8,     0, "::B:::::B:::W:W:"),
	(0,     0,     1,     ':',     14,     0, "::B:::::B:::W:W:"),
	(0,     0,     1,     'B',     11,     0, "::B:::::B:::W:W:"),
	(0,     0,     0,     'B',     7,     0, "::B:::::B::BW:W:"),
	(0,     1,     1,     'B',     14,     0, "::B:::::B::BW:W:"),
	(0,     0,     1,     'W',     10,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     7,     0, "::::::::::W:::B:"),
	(0,     0,     0,     ':',     8,     0, ":::::::W::W:::B:"),
	(0,     0,     1,     '*',     4,     0, ":::::::W::W:::B:"),
	(0,     0,     1,     'B',     11,     0, "::::*::W::W:::B:"),
	(0,     0,     0,     '*',     6,     0, "::::*::W::WB::B:"),
	(0,     0,     1,     '*',     15,     0, "::::*::W::WB::B:"),
	(0,     0,     1,     '*',     10,     0, "::::*::W::WB::B*"),
	(0,     0,     0,     ':',     12,     0, "::::*::W::BB::B*"),
	(0,     0,     1,     ':',     14,     0, "::::*::W::BB::B*"),
	(0,     0,     0,     ':',     13,     0, "::::*::W::BB::B*"),
	(0,     0,     0,     ':',     9,     0, "::::*::W::BB::B*"),
	(0,     1,     1,     'W',     12,     0, "::::*::W::BB::B*"),
	(0,     0,     0,     ':',     11,     0, "::::::::::::W:::"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::W:::"),
	(0,     0,     0,     'B',     7,     0, "::::::::::::W:::"),
	(0,     0,     1,     ':',     1,     0, "::::::::::::W:::"),
	(0,     0,     1,     'B',     3,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     10,     0, ":::B::::::::W:::"),
	(0,     0,     0,     'B',     15,     0, ":::B::::::::W:::"),
	(0,     0,     1,     '*',     1,     0, ":::B::::::::W:::"),
	(0,     1,     0,     ':',     14,     0, ":*:B::::::::W:::"),
	(0,     0,     0,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     15,     0, ":::::::::W::::::"),
	(0,     0,     0,     '*',     4,     0, ":::::::::W::::::"),
	(0,     0,     0,     'W',     11,     0, ":::::::::W::::::"),
	(0,     0,     1,     ':',     3,     0, ":::::::::W::::::"),
	(0,     0,     0,     'B',     10,     0, ":::::::::W::::::"),
	(0,     0,     0,     'B',     3,     0, ":::::::::W::::::"),
	(0,     1,     0,     'B',     5,     0, ":::::::::W::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::::::::::::W:"),
	(0,     0,     0,     'W',     14,     0, "::::::::::::::W:"),
	(0,     0,     1,     'W',     11,     0, "::::::::::::::W:"),
	(0,     0,     1,     '*',     2,     0, ":::::::::::W::W:"),
	(0,     0,     1,     'W',     7,     0, "::*::::::::W::W:"),
	(0,     0,     0,     '*',     4,     0, "::*::::W:::W::W:"),
	(0,     0,     0,     '*',     5,     0, "::*::::W:::W::W:"),
	(0,     0,     1,     'W',     7,     0, "::*::::W:::W::W:"),
	(0,     0,     0,     ':',     13,     0, "::*::::W:::W::W:"),
	(0,     0,     0,     ':',     12,     0, "::*::::W:::W::W:"),
	(0,     0,     0,     ':',     7,     0, "::*::::W:::W::W:"),
	(0,     0,     0,     'B',     1,     0, "::*::::W:::W::W:"),
	(0,     0,     1,     ':',     12,     0, "::*::::W:::W::W:"),
	(0,     0,     1,     'B',     7,     0, "::*::::W:::W::W:"),
	(0,     0,     1,     'B',     3,     0, "::*::::B:::W::W:"),
	(0,     0,     0,     '*',     8,     0, "::*B:::B:::W::W:"),
	(0,     1,     1,     'B',     6,     0, "::*B:::B:::W::W:"),
	(0,     0,     0,     'B',     1,     0, "::::::B:::::::::"),
	(0,     0,     0,     'W',     9,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     4,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::B:::::::::"),
	(0,     0,     1,     'W',     11,     0, "::::::B:::::::::"),
	(0,     1,     1,     'W',     6,     0, "::::::B::::W::::"),
	(0,     0,     0,     'B',     1,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     8,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     8,     0, "::::::W:B:::::::"),
	(0,     0,     1,     'W',     1,     0, "::::::W:B:::::::"),
	(0,     1,     1,     ':',     5,     0, ":W::::W:B:::::::"),
	(0,     1,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     0, ":::::B::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::::B::::::::::"),
	(0,     0,     0,     'W',     11,     0, ":::::B::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::B::::::::::"),
	(0,     0,     0,     ':',     10,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     12,     0, ":::::B::::::::::"),
	(0,     0,     0,     '*',     1,     0, ":::::B::::::B:::"),
	(0,     0,     0,     'B',     8,     0, ":::::B::::::B:::"),
	(0,     0,     0,     '*',     9,     0, ":::::B::::::B:::"),
	(0,     0,     1,     'W',     15,     0, ":::::B::::::B:::"),
	(0,     0,     1,     'W',     14,     0, ":::::B::::::B::W"),
	(0,     0,     0,     'B',     9,     0, ":::::B::::::B:WW"),
	(0,     0,     1,     '*',     3,     0, ":::::B::::::B:WW"),
	(0,     0,     0,     '*',     7,     0, ":::*:B::::::B:WW"),
	(0,     0,     0,     'W',     2,     0, ":::*:B::::::B:WW"),
	(0,     0,     1,     'B',     15,     0, ":::*:B::::::B:WW"),
	(0,     0,     0,     'B',     2,     0, ":::*:B::::::B:WB"),
	(0,     0,     0,     'W',     13,     0, ":::*:B::::::B:WB"),
	(0,     0,     1,     ':',     9,     0, ":::*:B::::::B:WB"),
	(0,     1,     0,     'W',     11,     0, ":::*:B::::::B:WB"),
	(0,     1,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     14,     0, ":::::W::::::::::"),
	(0,     1,     0,     'B',     13,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":::::::::W::::::"),
	(0,     0,     0,     ':',     7,     0, ":::::::::W:::*::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::W:::*::"),
	(0,     0,     0,     'B',     4,     0, ":::::::::W:::*::"),
	(0,     0,     1,     'B',     5,     0, ":::::::::W:::*::"),
	(0,     0,     1,     ':',     10,     0, ":::::B:::W:::*::"),
	(0,     0,     0,     ':',     4,     0, ":::::B:::W:::*::"),
	(0,     0,     1,     'B',     2,     0, ":::::B:::W:::*::"),
	(0,     0,     1,     '*',     13,     0, "::B::B:::W:::*::"),
	(0,     0,     1,     'W',     8,     0, "::B::B:::W::::::"),
	(0,     0,     0,     '*',     11,     0, "::B::B::WW::::::"),
	(0,     0,     1,     ':',     3,     0, "::B::B::WW::::::"),
	(0,     0,     0,     'B',     8,     0, "::B::B::WW::::::"),
	(0,     0,     1,     '*',     1,     0, "::B::B::WW::::::"),
	(0,     0,     0,     ':',     5,     0, ":*B::B::WW::::::"),
	(0,     0,     1,     '*',     1,     0, ":*B::B::WW::::::"),
	(0,     0,     0,     ':',     15,     0, "::B::B::WW::::::"),
	(0,     0,     0,     '*',     6,     0, "::B::B::WW::::::"),
	(0,     0,     1,     ':',     1,     0, "::B::B::WW::::::"),
	(0,     0,     0,     ':',     8,     0, "::B::B::WW::::::"),
	(0,     1,     0,     '*',     13,     0, "::B::B::WW::::::"),
	(0,     0,     0,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     5,     0, "::::::::::::::*:"),
	(0,     0,     1,     'B',     2,     0, "::::::::::::::*:"),
	(0,     0,     0,     '*',     12,     0, "::B:::::::::::*:"),
	(0,     1,     0,     'B',     7,     0, "::B:::::::::::*:"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     0, "W:::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "W:::::W:::::::::"),
	(0,     0,     0,     'B',     10,     0, "W:::W:W:::::::::"),
	(0,     0,     1,     '*',     8,     0, "W:::W:W:::::::::"),
	(0,     0,     1,     ':',     13,     0, "W:::W:W:*:::::::"),
	(0,     0,     1,     '*',     8,     0, "W:::W:W:*:::::::"),
	(0,     1,     0,     'B',     12,     0, "W:::W:W:::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::::::::::::*:"),
	(0,     0,     0,     ':',     4,     0, "::::::::::::::*:"),
	(0,     0,     0,     '*',     6,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     8,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     10,     0, "::::::::::::::*:"),
	(0,     0,     1,     ':',     14,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     5,     0, "::::::::::::::*:"),
	(0,     0,     0,     ':',     8,     0, "::::::::::::::*:"),
	(0,     0,     1,     ':',     7,     0, "::::::::::::::*:"),
	(0,     0,     0,     'B',     10,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     0,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     3,     0, "*:::::::::::::*:"),
	(0,     0,     1,     '*',     6,     0, "*:::::::::::::*:"),
	(0,     0,     0,     'B',     7,     0, "*:::::*:::::::*:"),
	(0,     0,     0,     ':',     3,     0, "*:::::*:::::::*:"),
	(0,     0,     1,     ':',     0,     0, "*:::::*:::::::*:"),
	(0,     0,     1,     '*',     2,     0, "*:::::*:::::::*:"),
	(0,     0,     1,     'W',     13,     0, "*:*:::*:::::::*:"),
	(0,     0,     1,     '*',     4,     0, "*:*:::*::::::W*:"),
	(0,     0,     1,     ':',     5,     0, "*:*:*:*::::::W*:"),
	(0,     0,     1,     ':',     7,     0, "*:*:*:*::::::W*:"),
	(0,     0,     1,     'B',     15,     0, "*:*:*:*::::::W*:"),
	(0,     0,     0,     ':',     1,     0, "*:*:*:*::::::W*B"),
	(0,     0,     0,     'W',     15,     0, "*:*:*:*::::::W*B"),
	(0,     0,     0,     'W',     3,     0, "*:*:*:*::::::W*B"),
	(0,     0,     1,     'B',     7,     0, "*:*:*:*::::::W*B"),
	(0,     0,     0,     'W',     14,     0, "*:*:*:*B:::::W*B"),
	(0,     1,     0,     'B',     8,     0, "*:*:*:*B:::::W*B"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     10,     0, ":::::B::::::::::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     0, "::B:::::::::::::"),
	(0,     1,     0,     'B',     3,     0, "::B:::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     8,     0, "::::::::::::::*:"),
	(0,     0,     0,     ':',     7,     0, "::::::::*:::::*:"),
	(0,     0,     0,     'B',     11,     0, "::::::::*:::::*:"),
	(0,     1,     0,     'W',     4,     0, "::::::::*:::::*:"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     9,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     9,     0, ":::*::::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::*::::::::::::"),
	(0,     0,     1,     'B',     9,     0, ":::*::::::::::::"),
	(0,     0,     0,     ':',     10,     0, ":::*:::::B::::::"),
	(0,     0,     1,     '*',     6,     0, ":::*:::::B::::::"),
	(0,     0,     1,     'W',     14,     0, ":::*::*::B::::::"),
	(0,     0,     0,     '*',     1,     0, ":::*::*::B::::W:"),
	(0,     0,     1,     '*',     8,     0, ":::*::*::B::::W:"),
	(0,     0,     1,     'B',     5,     0, ":::*::*:*B::::W:"),
	(0,     0,     0,     ':',     12,     0, ":::*:B*:*B::::W:"),
	(0,     0,     0,     '*',     11,     0, ":::*:B*:*B::::W:"),
	(0,     0,     0,     '*',     3,     0, ":::*:B*:*B::::W:"),
	(0,     0,     1,     '*',     11,     0, ":::*:B*:*B::::W:"),
	(0,     0,     1,     ':',     12,     0, ":::*:B*:*B:*::W:"),
	(0,     0,     1,     'B',     10,     0, ":::*:B*:*B:*::W:"),
	(0,     0,     1,     'B',     1,     0, ":::*:B*:*BB*::W:"),
	(0,     0,     1,     '*',     7,     0, ":B:*:B*:*BB*::W:"),
	(0,     0,     1,     'B',     8,     0, ":B:*:B***BB*::W:"),
	(0,     0,     0,     'B',     1,     0, ":B:*:B**BBB*::W:"),
	(0,     0,     0,     '*',     9,     0, ":B:*:B**BBB*::W:"),
	(0,     0,     1,     ':',     14,     0, ":B:*:B**BBB*::W:"),
	(0,     0,     1,     'W',     11,     0, ":B:*:B**BBB*::W:"),
	(0,     0,     0,     'W',     12,     0, ":B:*:B**BBBW::W:"),
	(0,     0,     1,     'B',     0,     0, ":B:*:B**BBBW::W:"),
	(0,     0,     0,     ':',     10,     0, "BB:*:B**BBBW::W:"),
	(0,     0,     1,     'W',     11,     0, "BB:*:B**BBBW::W:"),
	(0,     1,     0,     ':',     12,     0, "BB:*:B**BBBW::W:"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     0, ":::::::*::::::::"),
	(0,     0,     0,     '*',     7,     0, "::*::::*::::::::"),
	(0,     0,     1,     '*',     12,     0, "::*::::*::::::::"),
	(0,     0,     0,     ':',     8,     0, "::*::::*::::*:::"),
	(0,     0,     1,     'W',     3,     0, "::*::::*::::*:::"),
	(0,     0,     1,     '*',     8,     0, "::*W:::*::::*:::"),
	(0,     0,     1,     'B',     2,     0, "::*W:::**:::*:::"),
	(0,     0,     0,     ':',     13,     0, "::BW:::**:::*:::"),
	(0,     1,     1,     'B',     6,     0, "::BW:::**:::*:::"),
	(0,     0,     0,     'W',     14,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     14,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     1,     0, "::::::B:::::::::"),
	(0,     0,     1,     'B',     8,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     3,     0, "::::::B:B:::::::"),
	(0,     0,     1,     'B',     12,     0, "::::::B:B:::::::"),
	(0,     0,     0,     '*',     6,     0, "::::::B:B:::B:::"),
	(0,     1,     0,     ':',     15,     0, "::::::B:B:::B:::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     9,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::W:::::::::"),
	(0,     0,     0,     '*',     5,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     6,     0, "::::::W:::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     1,     0, "::*:::W:::::::::"),
	(0,     0,     0,     'B',     2,     0, ":B*:::W:::::::::"),
	(0,     0,     0,     'B',     13,     0, ":B*:::W:::::::::"),
	(0,     0,     1,     'W',     4,     0, ":B*:::W:::::::::"),
	(0,     0,     0,     ':',     14,     0, ":B*:W:W:::::::::")
	);
END PACKAGE ex4_data_pak;
